NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.01 ;

DIVIDERCHAR "/" ;
#MINFEATURE 0.001 0.001 ;


#LAYER GRLOGIC
#  TYPE  MASTERSLICE ;
#END GRLOGIC

#LAYER NW
#  TYPE	MASTERSLICE ;
#END NW

#LAYER RX
#  TYPE	MASTERSLICE ;
#END RX

#LAYER BP
#  TYPE	MASTERSLICE ;
#END BP

#LAYER PC
#  TYPE	MASTERSLICE ;
#END PC

#LAYER CA
#  TYPE	CUT ;
#END CA

LAYER M1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		CUSTOM_PITCH ;
  WIDTH		0.16 ;
  AREA		0.12 ;
  SPACING	0.16 ;
  SPACING	0.26 RANGE 1.76 4 ;
  SPACING	0.36 RANGE 4 8 ;
  SPACING	1.12 RANGE 8 25 ;
  SPACING	1.92 RANGE 25 100000 ;
END M1

LAYER V1
  TYPE	CUT ;
END V1

LAYER M2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		CUSTOM_PITCH ;
  WIDTH		0.2 ;
  AREA		0.12 ;
  SPACING	0.2 ;
  SPACING	0.28 RANGE 2 4 ;
  SPACING	0.36 RANGE 4 8 ;
  SPACING	1.12 RANGE 8 25 ;
  SPACING	1.92 RANGE 25 100000 ;
  CURRENTDEN 0 ;
END M2

LAYER V2
  TYPE	CUT ;
END V2

LAYER M3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		CUSTOM_PITCH ;
  WIDTH		0.2 ;
  AREA		0.12 ;
  SPACING	0.2 ;
  SPACING	0.28 RANGE 2 4 ;
  SPACING	0.36 RANGE 4 8 ;
  SPACING	1.12 RANGE 8 25 ;
  SPACING	1.92 RANGE 25 100000 ;
END M3

LAYER V3
  TYPE	CUT ;
END V3

LAYER M4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		CUSTOM_PITCH ;
  WIDTH		0.2 ;
  AREA		0.12 ;
  SPACING	0.2 ;
  SPACING	0.28 RANGE 2 4 ;
  SPACING	0.36 RANGE 4 8 ;
  SPACING	1.12 RANGE 8 25 ;
  SPACING	1.92 RANGE 25 100000 ;
END M4

LAYER V4
  TYPE	CUT ;
END V4

LAYER M5
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		CUSTOM_PITCH ;
  WIDTH		0.2 ;
  AREA		0.12 ;
  SPACING	0.2 ;
  SPACING	0.28 RANGE 2 4 ;
  SPACING	0.36 RANGE 4 8 ;
  SPACING	1.12 RANGE 8 25 ;
  SPACING	1.92 RANGE 25 100000 ;
END M5

LAYER V5
  TYPE	CUT ;
END V5

LAYER M6
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		CUSTOM_PITCH ;
  WIDTH		0.2 ;
  AREA		0.12 ;
  SPACING	0.2 ;
  SPACING	0.28 RANGE 2 4 ;
  SPACING	0.36 RANGE 4 8 ;
  SPACING	1.12 RANGE 8 25 ;
  SPACING	1.92 RANGE 25 100000 ;
END M6

LAYER OVERLAP
  TYPE	OVERLAP ;
END OVERLAP

SPACING
  SAMENET M1  M1	0.16 STACK ;
  SAMENET M2  M2	0.2 STACK ;
  SAMENET M3  M3	0.2 STACK ;
  SAMENET M4  M4	0.2 STACK ;
  SAMENET M5  M5	0.2 STACK ;
  SAMENET M6  M6	0.2 STACK ;
  SAMENET V1  V1	0.2 ;
  SAMENET V2  V2	0.2 ;
  SAMENET V3  V3	0.2 ;
  SAMENET V4  V4	0.2 ;
  SAMENET V5  V5	0.2 ;
  SAMENET V1  V2	0.00 STACK ;
  SAMENET V2  V3	0.00 STACK ;
  SAMENET V3  V4	0.00 STACK ;
  SAMENET V4  V5	0.00 STACK ;
  SAMENET V1  V3	0.00 STACK ;
  SAMENET V2  V4	0.00 STACK ;
  SAMENET V3  V5	0.00 STACK ;
  SAMENET V1  V4	0.00 STACK ;
  SAMENET V2  V5	0.00 STACK ;
  SAMENET V1  V5	0.00 STACK ;
END SPACING

VIA via5 DEFAULT
  LAYER M5 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER V5 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER M6 ;
    RECT -0.1 -0.1 0.1 0.1 ;
END via5

VIA via4 DEFAULT
  LAYER M4 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER V4 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER M5 ;
    RECT -0.1 -0.1 0.1 0.1 ;
END via4

VIA via3 DEFAULT
  LAYER M4 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER V3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER M3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
END via3

VIA via2 DEFAULT
  LAYER M3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER V2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER M2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
END via2

VIA via1 DEFAULT
  LAYER M2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER V1 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER M1 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END via1

VIARULE via1Array GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.09 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.09 ;
    METALOVERHANG 0 ;
  LAYER V1 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
END via1Array

VIARULE via2Array GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER V2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
END via2Array

VIARULE via3Array GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER V3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
END via3Array

VIARULE via4Array GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER V4 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
END via4Array

VIARULE via5Array GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.09 ;
    METALOVERHANG 0 ;
  LAYER V5 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
END via5Array

VIARULE TURNM1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
  LAYER M1 ;
    DIRECTION VERTICAL ;
END TURNM1

VIARULE TURNM2 GENERATE
  LAYER M2 ;
    DIRECTION HORIZONTAL ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
END TURNM2

VIARULE TURNM3 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
  LAYER M3 ;
    DIRECTION VERTICAL ;
END TURNM3

VIARULE TURNM4 GENERATE
  LAYER M4 ;
    DIRECTION HORIZONTAL ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
END TURNM4

VIARULE TURNM5 GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
  LAYER M5 ;
    DIRECTION VERTICAL ;
END TURNM5

VIARULE TURNM6 GENERATE
  LAYER M6 ;
    DIRECTION HORIZONTAL ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
END TURNM6

