module inv(a, out);
input a;
output out;
assign out = ~a;
endmodule

module nand2(a, b, out);
input a, b;
output out;
assign out = ~(a & b);
endmodule

module xor2(a, b, out);
input a, b;
output out;
assign out = (a ^ b);
endmodule

module d_ff( D, clk, R, Q);
input D, clk, R;
output Q;
reg Q;
always @(posedge clk or negedge R)
  if (R == 1'b1)
    Q = 1'b0;
  else
    Q = D;
endmodule


/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : L-2016.03-SP3
// Date      : Mon Sep 24 07:58:36 2018
/////////////////////////////////////////////////////////////


module decoder1024 ( out, clk, clr, enable, sig, prgm );
  input clk, clr, enable, sig, prgm;
  output out;
  wire   \prgm_register/n2048 , \prgm_register/n2047 , \prgm_register/n2046 ,
         \prgm_register/n2045 , \prgm_register/n2044 , \prgm_register/n2043 ,
         \prgm_register/n2042 , \prgm_register/n2041 , \prgm_register/n2040 ,
         \prgm_register/n2039 , \prgm_register/n2038 , \prgm_register/n2037 ,
         \prgm_register/n2036 , \prgm_register/n2035 , \prgm_register/n2034 ,
         \prgm_register/n2033 , \prgm_register/n2032 , \prgm_register/n2031 ,
         \prgm_register/n2030 , \prgm_register/n2029 , \prgm_register/n2028 ,
         \prgm_register/n2027 , \prgm_register/n2026 , \prgm_register/n2025 ,
         \prgm_register/n2024 , \prgm_register/n2023 , \prgm_register/n2022 ,
         \prgm_register/n2021 , \prgm_register/n2020 , \prgm_register/n2019 ,
         \prgm_register/n2018 , \prgm_register/n2017 , \prgm_register/n2016 ,
         \prgm_register/n2015 , \prgm_register/n2014 , \prgm_register/n2013 ,
         \prgm_register/n2012 , \prgm_register/n2011 , \prgm_register/n2010 ,
         \prgm_register/n2009 , \prgm_register/n2008 , \prgm_register/n2007 ,
         \prgm_register/n2006 , \prgm_register/n2005 , \prgm_register/n2004 ,
         \prgm_register/n2003 , \prgm_register/n2002 , \prgm_register/n2001 ,
         \prgm_register/n2000 , \prgm_register/n1999 , \prgm_register/n1998 ,
         \prgm_register/n1997 , \prgm_register/n1996 , \prgm_register/n1995 ,
         \prgm_register/n1994 , \prgm_register/n1993 , \prgm_register/n1992 ,
         \prgm_register/n1991 , \prgm_register/n1990 , \prgm_register/n1989 ,
         \prgm_register/n1988 , \prgm_register/n1987 , \prgm_register/n1986 ,
         \prgm_register/n1985 , \prgm_register/n1984 , \prgm_register/n1983 ,
         \prgm_register/n1982 , \prgm_register/n1981 , \prgm_register/n1980 ,
         \prgm_register/n1979 , \prgm_register/n1978 , \prgm_register/n1977 ,
         \prgm_register/n1976 , \prgm_register/n1975 , \prgm_register/n1974 ,
         \prgm_register/n1973 , \prgm_register/n1972 , \prgm_register/n1971 ,
         \prgm_register/n1970 , \prgm_register/n1969 , \prgm_register/n1968 ,
         \prgm_register/n1967 , \prgm_register/n1966 , \prgm_register/n1965 ,
         \prgm_register/n1964 , \prgm_register/n1963 , \prgm_register/n1962 ,
         \prgm_register/n1961 , \prgm_register/n1960 , \prgm_register/n1959 ,
         \prgm_register/n1958 , \prgm_register/n1957 , \prgm_register/n1956 ,
         \prgm_register/n1955 , \prgm_register/n1954 , \prgm_register/n1953 ,
         \prgm_register/n1952 , \prgm_register/n1951 , \prgm_register/n1950 ,
         \prgm_register/n1949 , \prgm_register/n1948 , \prgm_register/n1947 ,
         \prgm_register/n1946 , \prgm_register/n1945 , \prgm_register/n1944 ,
         \prgm_register/n1943 , \prgm_register/n1942 , \prgm_register/n1941 ,
         \prgm_register/n1940 , \prgm_register/n1939 , \prgm_register/n1938 ,
         \prgm_register/n1937 , \prgm_register/n1936 , \prgm_register/n1935 ,
         \prgm_register/n1934 , \prgm_register/n1933 , \prgm_register/n1932 ,
         \prgm_register/n1931 , \prgm_register/n1930 , \prgm_register/n1929 ,
         \prgm_register/n1928 , \prgm_register/n1927 , \prgm_register/n1926 ,
         \prgm_register/n1925 , \prgm_register/n1924 , \prgm_register/n1923 ,
         \prgm_register/n1922 , \prgm_register/n1921 , \prgm_register/n1920 ,
         \prgm_register/n1919 , \prgm_register/n1918 , \prgm_register/n1917 ,
         \prgm_register/n1916 , \prgm_register/n1915 , \prgm_register/n1914 ,
         \prgm_register/n1913 , \prgm_register/n1912 , \prgm_register/n1911 ,
         \prgm_register/n1910 , \prgm_register/n1909 , \prgm_register/n1908 ,
         \prgm_register/n1907 , \prgm_register/n1906 , \prgm_register/n1905 ,
         \prgm_register/n1904 , \prgm_register/n1903 , \prgm_register/n1902 ,
         \prgm_register/n1901 , \prgm_register/n1900 , \prgm_register/n1899 ,
         \prgm_register/n1898 , \prgm_register/n1897 , \prgm_register/n1896 ,
         \prgm_register/n1895 , \prgm_register/n1894 , \prgm_register/n1893 ,
         \prgm_register/n1892 , \prgm_register/n1891 , \prgm_register/n1890 ,
         \prgm_register/n1889 , \prgm_register/n1888 , \prgm_register/n1887 ,
         \prgm_register/n1886 , \prgm_register/n1885 , \prgm_register/n1884 ,
         \prgm_register/n1883 , \prgm_register/n1882 , \prgm_register/n1881 ,
         \prgm_register/n1880 , \prgm_register/n1879 , \prgm_register/n1878 ,
         \prgm_register/n1877 , \prgm_register/n1876 , \prgm_register/n1875 ,
         \prgm_register/n1874 , \prgm_register/n1873 , \prgm_register/n1872 ,
         \prgm_register/n1871 , \prgm_register/n1870 , \prgm_register/n1869 ,
         \prgm_register/n1868 , \prgm_register/n1867 , \prgm_register/n1866 ,
         \prgm_register/n1865 , \prgm_register/n1864 , \prgm_register/n1863 ,
         \prgm_register/n1862 , \prgm_register/n1861 , \prgm_register/n1860 ,
         \prgm_register/n1859 , \prgm_register/n1858 , \prgm_register/n1857 ,
         \prgm_register/n1856 , \prgm_register/n1855 , \prgm_register/n1854 ,
         \prgm_register/n1853 , \prgm_register/n1852 , \prgm_register/n1851 ,
         \prgm_register/n1850 , \prgm_register/n1849 , \prgm_register/n1848 ,
         \prgm_register/n1847 , \prgm_register/n1846 , \prgm_register/n1845 ,
         \prgm_register/n1844 , \prgm_register/n1843 , \prgm_register/n1842 ,
         \prgm_register/n1841 , \prgm_register/n1840 , \prgm_register/n1839 ,
         \prgm_register/n1838 , \prgm_register/n1837 , \prgm_register/n1836 ,
         \prgm_register/n1835 , \prgm_register/n1834 , \prgm_register/n1833 ,
         \prgm_register/n1832 , \prgm_register/n1831 , \prgm_register/n1830 ,
         \prgm_register/n1829 , \prgm_register/n1828 , \prgm_register/n1827 ,
         \prgm_register/n1826 , \prgm_register/n1825 , \prgm_register/n1824 ,
         \prgm_register/n1823 , \prgm_register/n1822 , \prgm_register/n1821 ,
         \prgm_register/n1820 , \prgm_register/n1819 , \prgm_register/n1818 ,
         \prgm_register/n1817 , \prgm_register/n1816 , \prgm_register/n1815 ,
         \prgm_register/n1814 , \prgm_register/n1813 , \prgm_register/n1812 ,
         \prgm_register/n1811 , \prgm_register/n1810 , \prgm_register/n1809 ,
         \prgm_register/n1808 , \prgm_register/n1807 , \prgm_register/n1806 ,
         \prgm_register/n1805 , \prgm_register/n1804 , \prgm_register/n1803 ,
         \prgm_register/n1802 , \prgm_register/n1801 , \prgm_register/n1800 ,
         \prgm_register/n1799 , \prgm_register/n1798 , \prgm_register/n1797 ,
         \prgm_register/n1796 , \prgm_register/n1795 , \prgm_register/n1794 ,
         \prgm_register/n1793 , \prgm_register/n1792 , \prgm_register/n1791 ,
         \prgm_register/n1790 , \prgm_register/n1789 , \prgm_register/n1788 ,
         \prgm_register/n1787 , \prgm_register/n1786 , \prgm_register/n1785 ,
         \prgm_register/n1784 , \prgm_register/n1783 , \prgm_register/n1782 ,
         \prgm_register/n1781 , \prgm_register/n1780 , \prgm_register/n1779 ,
         \prgm_register/n1778 , \prgm_register/n1777 , \prgm_register/n1776 ,
         \prgm_register/n1775 , \prgm_register/n1774 , \prgm_register/n1773 ,
         \prgm_register/n1772 , \prgm_register/n1771 , \prgm_register/n1770 ,
         \prgm_register/n1769 , \prgm_register/n1768 , \prgm_register/n1767 ,
         \prgm_register/n1766 , \prgm_register/n1765 , \prgm_register/n1764 ,
         \prgm_register/n1763 , \prgm_register/n1762 , \prgm_register/n1761 ,
         \prgm_register/n1760 , \prgm_register/n1759 , \prgm_register/n1758 ,
         \prgm_register/n1757 , \prgm_register/n1756 , \prgm_register/n1755 ,
         \prgm_register/n1754 , \prgm_register/n1753 , \prgm_register/n1752 ,
         \prgm_register/n1751 , \prgm_register/n1750 , \prgm_register/n1749 ,
         \prgm_register/n1748 , \prgm_register/n1747 , \prgm_register/n1746 ,
         \prgm_register/n1745 , \prgm_register/n1744 , \prgm_register/n1743 ,
         \prgm_register/n1742 , \prgm_register/n1741 , \prgm_register/n1740 ,
         \prgm_register/n1739 , \prgm_register/n1738 , \prgm_register/n1737 ,
         \prgm_register/n1736 , \prgm_register/n1735 , \prgm_register/n1734 ,
         \prgm_register/n1733 , \prgm_register/n1732 , \prgm_register/n1731 ,
         \prgm_register/n1730 , \prgm_register/n1729 , \prgm_register/n1728 ,
         \prgm_register/n1727 , \prgm_register/n1726 , \prgm_register/n1725 ,
         \prgm_register/n1724 , \prgm_register/n1723 , \prgm_register/n1722 ,
         \prgm_register/n1721 , \prgm_register/n1720 , \prgm_register/n1719 ,
         \prgm_register/n1718 , \prgm_register/n1717 , \prgm_register/n1716 ,
         \prgm_register/n1715 , \prgm_register/n1714 , \prgm_register/n1713 ,
         \prgm_register/n1712 , \prgm_register/n1711 , \prgm_register/n1710 ,
         \prgm_register/n1709 , \prgm_register/n1708 , \prgm_register/n1707 ,
         \prgm_register/n1706 , \prgm_register/n1705 , \prgm_register/n1704 ,
         \prgm_register/n1703 , \prgm_register/n1702 , \prgm_register/n1701 ,
         \prgm_register/n1700 , \prgm_register/n1699 , \prgm_register/n1698 ,
         \prgm_register/n1697 , \prgm_register/n1696 , \prgm_register/n1695 ,
         \prgm_register/n1694 , \prgm_register/n1693 , \prgm_register/n1692 ,
         \prgm_register/n1691 , \prgm_register/n1690 , \prgm_register/n1689 ,
         \prgm_register/n1688 , \prgm_register/n1687 , \prgm_register/n1686 ,
         \prgm_register/n1685 , \prgm_register/n1684 , \prgm_register/n1683 ,
         \prgm_register/n1682 , \prgm_register/n1681 , \prgm_register/n1680 ,
         \prgm_register/n1679 , \prgm_register/n1678 , \prgm_register/n1677 ,
         \prgm_register/n1676 , \prgm_register/n1675 , \prgm_register/n1674 ,
         \prgm_register/n1673 , \prgm_register/n1672 , \prgm_register/n1671 ,
         \prgm_register/n1670 , \prgm_register/n1669 , \prgm_register/n1668 ,
         \prgm_register/n1667 , \prgm_register/n1666 , \prgm_register/n1665 ,
         \prgm_register/n1664 , \prgm_register/n1663 , \prgm_register/n1662 ,
         \prgm_register/n1661 , \prgm_register/n1660 , \prgm_register/n1659 ,
         \prgm_register/n1658 , \prgm_register/n1657 , \prgm_register/n1656 ,
         \prgm_register/n1655 , \prgm_register/n1654 , \prgm_register/n1653 ,
         \prgm_register/n1652 , \prgm_register/n1651 , \prgm_register/n1650 ,
         \prgm_register/n1649 , \prgm_register/n1648 , \prgm_register/n1647 ,
         \prgm_register/n1646 , \prgm_register/n1645 , \prgm_register/n1644 ,
         \prgm_register/n1643 , \prgm_register/n1642 , \prgm_register/n1641 ,
         \prgm_register/n1640 , \prgm_register/n1639 , \prgm_register/n1638 ,
         \prgm_register/n1637 , \prgm_register/n1636 , \prgm_register/n1635 ,
         \prgm_register/n1634 , \prgm_register/n1633 , \prgm_register/n1632 ,
         \prgm_register/n1631 , \prgm_register/n1630 , \prgm_register/n1629 ,
         \prgm_register/n1628 , \prgm_register/n1627 , \prgm_register/n1626 ,
         \prgm_register/n1625 , \prgm_register/n1624 , \prgm_register/n1623 ,
         \prgm_register/n1622 , \prgm_register/n1621 , \prgm_register/n1620 ,
         \prgm_register/n1619 , \prgm_register/n1618 , \prgm_register/n1617 ,
         \prgm_register/n1616 , \prgm_register/n1615 , \prgm_register/n1614 ,
         \prgm_register/n1613 , \prgm_register/n1612 , \prgm_register/n1611 ,
         \prgm_register/n1610 , \prgm_register/n1609 , \prgm_register/n1608 ,
         \prgm_register/n1607 , \prgm_register/n1606 , \prgm_register/n1605 ,
         \prgm_register/n1604 , \prgm_register/n1603 , \prgm_register/n1602 ,
         \prgm_register/n1601 , \prgm_register/n1600 , \prgm_register/n1599 ,
         \prgm_register/n1598 , \prgm_register/n1597 , \prgm_register/n1596 ,
         \prgm_register/n1595 , \prgm_register/n1594 , \prgm_register/n1593 ,
         \prgm_register/n1592 , \prgm_register/n1591 , \prgm_register/n1590 ,
         \prgm_register/n1589 , \prgm_register/n1588 , \prgm_register/n1587 ,
         \prgm_register/n1586 , \prgm_register/n1585 , \prgm_register/n1584 ,
         \prgm_register/n1583 , \prgm_register/n1582 , \prgm_register/n1581 ,
         \prgm_register/n1580 , \prgm_register/n1579 , \prgm_register/n1578 ,
         \prgm_register/n1577 , \prgm_register/n1576 , \prgm_register/n1575 ,
         \prgm_register/n1574 , \prgm_register/n1573 , \prgm_register/n1572 ,
         \prgm_register/n1571 , \prgm_register/n1570 , \prgm_register/n1569 ,
         \prgm_register/n1568 , \prgm_register/n1567 , \prgm_register/n1566 ,
         \prgm_register/n1565 , \prgm_register/n1564 , \prgm_register/n1563 ,
         \prgm_register/n1562 , \prgm_register/n1561 , \prgm_register/n1560 ,
         \prgm_register/n1559 , \prgm_register/n1558 , \prgm_register/n1557 ,
         \prgm_register/n1556 , \prgm_register/n1555 , \prgm_register/n1554 ,
         \prgm_register/n1553 , \prgm_register/n1552 , \prgm_register/n1551 ,
         \prgm_register/n1550 , \prgm_register/n1549 , \prgm_register/n1548 ,
         \prgm_register/n1547 , \prgm_register/n1546 , \prgm_register/n1545 ,
         \prgm_register/n1544 , \prgm_register/n1543 , \prgm_register/n1542 ,
         \prgm_register/n1541 , \prgm_register/n1540 , \prgm_register/n1539 ,
         \prgm_register/n1538 , \prgm_register/n1537 , \prgm_register/n1536 ,
         \prgm_register/n1535 , \prgm_register/n1534 , \prgm_register/n1533 ,
         \prgm_register/n1532 , \prgm_register/n1531 , \prgm_register/n1530 ,
         \prgm_register/n1529 , \prgm_register/n1528 , \prgm_register/n1527 ,
         \prgm_register/n1526 , \prgm_register/n1525 , \prgm_register/n1524 ,
         \prgm_register/n1523 , \prgm_register/n1522 , \prgm_register/n1521 ,
         \prgm_register/n1520 , \prgm_register/n1519 , \prgm_register/n1518 ,
         \prgm_register/n1517 , \prgm_register/n1516 , \prgm_register/n1515 ,
         \prgm_register/n1514 , \prgm_register/n1513 , \prgm_register/n1512 ,
         \prgm_register/n1511 , \prgm_register/n1510 , \prgm_register/n1509 ,
         \prgm_register/n1508 , \prgm_register/n1507 , \prgm_register/n1506 ,
         \prgm_register/n1505 , \prgm_register/n1504 , \prgm_register/n1503 ,
         \prgm_register/n1502 , \prgm_register/n1501 , \prgm_register/n1500 ,
         \prgm_register/n1499 , \prgm_register/n1498 , \prgm_register/n1497 ,
         \prgm_register/n1496 , \prgm_register/n1495 , \prgm_register/n1494 ,
         \prgm_register/n1493 , \prgm_register/n1492 , \prgm_register/n1491 ,
         \prgm_register/n1490 , \prgm_register/n1489 , \prgm_register/n1488 ,
         \prgm_register/n1487 , \prgm_register/n1486 , \prgm_register/n1485 ,
         \prgm_register/n1484 , \prgm_register/n1483 , \prgm_register/n1482 ,
         \prgm_register/n1481 , \prgm_register/n1480 , \prgm_register/n1479 ,
         \prgm_register/n1478 , \prgm_register/n1477 , \prgm_register/n1476 ,
         \prgm_register/n1475 , \prgm_register/n1474 , \prgm_register/n1473 ,
         \prgm_register/n1472 , \prgm_register/n1471 , \prgm_register/n1470 ,
         \prgm_register/n1469 , \prgm_register/n1468 , \prgm_register/n1467 ,
         \prgm_register/n1466 , \prgm_register/n1465 , \prgm_register/n1464 ,
         \prgm_register/n1463 , \prgm_register/n1462 , \prgm_register/n1461 ,
         \prgm_register/n1460 , \prgm_register/n1459 , \prgm_register/n1458 ,
         \prgm_register/n1457 , \prgm_register/n1456 , \prgm_register/n1455 ,
         \prgm_register/n1454 , \prgm_register/n1453 , \prgm_register/n1452 ,
         \prgm_register/n1451 , \prgm_register/n1450 , \prgm_register/n1449 ,
         \prgm_register/n1448 , \prgm_register/n1447 , \prgm_register/n1446 ,
         \prgm_register/n1445 , \prgm_register/n1444 , \prgm_register/n1443 ,
         \prgm_register/n1442 , \prgm_register/n1441 , \prgm_register/n1440 ,
         \prgm_register/n1439 , \prgm_register/n1438 , \prgm_register/n1437 ,
         \prgm_register/n1436 , \prgm_register/n1435 , \prgm_register/n1434 ,
         \prgm_register/n1433 , \prgm_register/n1432 , \prgm_register/n1431 ,
         \prgm_register/n1430 , \prgm_register/n1429 , \prgm_register/n1428 ,
         \prgm_register/n1427 , \prgm_register/n1426 , \prgm_register/n1425 ,
         \prgm_register/n1424 , \prgm_register/n1423 , \prgm_register/n1422 ,
         \prgm_register/n1421 , \prgm_register/n1420 , \prgm_register/n1419 ,
         \prgm_register/n1418 , \prgm_register/n1417 , \prgm_register/n1416 ,
         \prgm_register/n1415 , \prgm_register/n1414 , \prgm_register/n1413 ,
         \prgm_register/n1412 , \prgm_register/n1411 , \prgm_register/n1410 ,
         \prgm_register/n1409 , \prgm_register/n1408 , \prgm_register/n1407 ,
         \prgm_register/n1406 , \prgm_register/n1405 , \prgm_register/n1404 ,
         \prgm_register/n1403 , \prgm_register/n1402 , \prgm_register/n1401 ,
         \prgm_register/n1400 , \prgm_register/n1399 , \prgm_register/n1398 ,
         \prgm_register/n1397 , \prgm_register/n1396 , \prgm_register/n1395 ,
         \prgm_register/n1394 , \prgm_register/n1393 , \prgm_register/n1392 ,
         \prgm_register/n1391 , \prgm_register/n1390 , \prgm_register/n1389 ,
         \prgm_register/n1388 , \prgm_register/n1387 , \prgm_register/n1386 ,
         \prgm_register/n1385 , \prgm_register/n1384 , \prgm_register/n1383 ,
         \prgm_register/n1382 , \prgm_register/n1381 , \prgm_register/n1380 ,
         \prgm_register/n1379 , \prgm_register/n1378 , \prgm_register/n1377 ,
         \prgm_register/n1376 , \prgm_register/n1375 , \prgm_register/n1374 ,
         \prgm_register/n1373 , \prgm_register/n1372 , \prgm_register/n1371 ,
         \prgm_register/n1370 , \prgm_register/n1369 , \prgm_register/n1368 ,
         \prgm_register/n1367 , \prgm_register/n1366 , \prgm_register/n1365 ,
         \prgm_register/n1364 , \prgm_register/n1363 , \prgm_register/n1362 ,
         \prgm_register/n1361 , \prgm_register/n1360 , \prgm_register/n1359 ,
         \prgm_register/n1358 , \prgm_register/n1357 , \prgm_register/n1356 ,
         \prgm_register/n1355 , \prgm_register/n1354 , \prgm_register/n1353 ,
         \prgm_register/n1352 , \prgm_register/n1351 , \prgm_register/n1350 ,
         \prgm_register/n1349 , \prgm_register/n1348 , \prgm_register/n1347 ,
         \prgm_register/n1346 , \prgm_register/n1345 , \prgm_register/n1344 ,
         \prgm_register/n1343 , \prgm_register/n1342 , \prgm_register/n1341 ,
         \prgm_register/n1340 , \prgm_register/n1339 , \prgm_register/n1338 ,
         \prgm_register/n1337 , \prgm_register/n1336 , \prgm_register/n1335 ,
         \prgm_register/n1334 , \prgm_register/n1333 , \prgm_register/n1332 ,
         \prgm_register/n1331 , \prgm_register/n1330 , \prgm_register/n1329 ,
         \prgm_register/n1328 , \prgm_register/n1327 , \prgm_register/n1326 ,
         \prgm_register/n1325 , \prgm_register/n1324 , \prgm_register/n1323 ,
         \prgm_register/n1322 , \prgm_register/n1321 , \prgm_register/n1320 ,
         \prgm_register/n1319 , \prgm_register/n1318 , \prgm_register/n1317 ,
         \prgm_register/n1316 , \prgm_register/n1315 , \prgm_register/n1314 ,
         \prgm_register/n1313 , \prgm_register/n1312 , \prgm_register/n1311 ,
         \prgm_register/n1310 , \prgm_register/n1309 , \prgm_register/n1308 ,
         \prgm_register/n1307 , \prgm_register/n1306 , \prgm_register/n1305 ,
         \prgm_register/n1304 , \prgm_register/n1303 , \prgm_register/n1302 ,
         \prgm_register/n1301 , \prgm_register/n1300 , \prgm_register/n1299 ,
         \prgm_register/n1298 , \prgm_register/n1297 , \prgm_register/n1296 ,
         \prgm_register/n1295 , \prgm_register/n1294 , \prgm_register/n1293 ,
         \prgm_register/n1292 , \prgm_register/n1291 , \prgm_register/n1290 ,
         \prgm_register/n1289 , \prgm_register/n1288 , \prgm_register/n1287 ,
         \prgm_register/n1286 , \prgm_register/n1285 , \prgm_register/n1284 ,
         \prgm_register/n1283 , \prgm_register/n1282 , \prgm_register/n1281 ,
         \prgm_register/n1280 , \prgm_register/n1279 , \prgm_register/n1278 ,
         \prgm_register/n1277 , \prgm_register/n1276 , \prgm_register/n1275 ,
         \prgm_register/n1274 , \prgm_register/n1273 , \prgm_register/n1272 ,
         \prgm_register/n1271 , \prgm_register/n1270 , \prgm_register/n1269 ,
         \prgm_register/n1268 , \prgm_register/n1267 , \prgm_register/n1266 ,
         \prgm_register/n1265 , \prgm_register/n1264 , \prgm_register/n1263 ,
         \prgm_register/n1262 , \prgm_register/n1261 , \prgm_register/n1260 ,
         \prgm_register/n1259 , \prgm_register/n1258 , \prgm_register/n1257 ,
         \prgm_register/n1256 , \prgm_register/n1255 , \prgm_register/n1254 ,
         \prgm_register/n1253 , \prgm_register/n1252 , \prgm_register/n1251 ,
         \prgm_register/n1250 , \prgm_register/n1249 , \prgm_register/n1248 ,
         \prgm_register/n1247 , \prgm_register/n1246 , \prgm_register/n1245 ,
         \prgm_register/n1244 , \prgm_register/n1243 , \prgm_register/n1242 ,
         \prgm_register/n1241 , \prgm_register/n1240 , \prgm_register/n1239 ,
         \prgm_register/n1238 , \prgm_register/n1237 , \prgm_register/n1236 ,
         \prgm_register/n1235 , \prgm_register/n1234 , \prgm_register/n1233 ,
         \prgm_register/n1232 , \prgm_register/n1231 , \prgm_register/n1230 ,
         \prgm_register/n1229 , \prgm_register/n1228 , \prgm_register/n1227 ,
         \prgm_register/n1226 , \prgm_register/n1225 , \prgm_register/n1224 ,
         \prgm_register/n1223 , \prgm_register/n1222 , \prgm_register/n1221 ,
         \prgm_register/n1220 , \prgm_register/n1219 , \prgm_register/n1218 ,
         \prgm_register/n1217 , \prgm_register/n1216 , \prgm_register/n1215 ,
         \prgm_register/n1214 , \prgm_register/n1213 , \prgm_register/n1212 ,
         \prgm_register/n1211 , \prgm_register/n1210 , \prgm_register/n1209 ,
         \prgm_register/n1208 , \prgm_register/n1207 , \prgm_register/n1206 ,
         \prgm_register/n1205 , \prgm_register/n1204 , \prgm_register/n1203 ,
         \prgm_register/n1202 , \prgm_register/n1201 , \prgm_register/n1200 ,
         \prgm_register/n1199 , \prgm_register/n1198 , \prgm_register/n1197 ,
         \prgm_register/n1196 , \prgm_register/n1195 , \prgm_register/n1194 ,
         \prgm_register/n1193 , \prgm_register/n1192 , \prgm_register/n1191 ,
         \prgm_register/n1190 , \prgm_register/n1189 , \prgm_register/n1188 ,
         \prgm_register/n1187 , \prgm_register/n1186 , \prgm_register/n1185 ,
         \prgm_register/n1184 , \prgm_register/n1183 , \prgm_register/n1182 ,
         \prgm_register/n1181 , \prgm_register/n1180 , \prgm_register/n1179 ,
         \prgm_register/n1178 , \prgm_register/n1177 , \prgm_register/n1176 ,
         \prgm_register/n1175 , \prgm_register/n1174 , \prgm_register/n1173 ,
         \prgm_register/n1172 , \prgm_register/n1171 , \prgm_register/n1170 ,
         \prgm_register/n1169 , \prgm_register/n1168 , \prgm_register/n1167 ,
         \prgm_register/n1166 , \prgm_register/n1165 , \prgm_register/n1164 ,
         \prgm_register/n1163 , \prgm_register/n1162 , \prgm_register/n1161 ,
         \prgm_register/n1160 , \prgm_register/n1159 , \prgm_register/n1158 ,
         \prgm_register/n1157 , \prgm_register/n1156 , \prgm_register/n1155 ,
         \prgm_register/n1154 , \prgm_register/n1153 , \prgm_register/n1152 ,
         \prgm_register/n1151 , \prgm_register/n1150 , \prgm_register/n1149 ,
         \prgm_register/n1148 , \prgm_register/n1147 , \prgm_register/n1146 ,
         \prgm_register/n1145 , \prgm_register/n1144 , \prgm_register/n1143 ,
         \prgm_register/n1142 , \prgm_register/n1141 , \prgm_register/n1140 ,
         \prgm_register/n1139 , \prgm_register/n1138 , \prgm_register/n1137 ,
         \prgm_register/n1136 , \prgm_register/n1135 , \prgm_register/n1134 ,
         \prgm_register/n1133 , \prgm_register/n1132 , \prgm_register/n1131 ,
         \prgm_register/n1130 , \prgm_register/n1129 , \prgm_register/n1128 ,
         \prgm_register/n1127 , \prgm_register/n1126 , \prgm_register/n1125 ,
         \prgm_register/n1124 , \prgm_register/n1123 , \prgm_register/n1122 ,
         \prgm_register/n1121 , \prgm_register/n1120 , \prgm_register/n1119 ,
         \prgm_register/n1118 , \prgm_register/n1117 , \prgm_register/n1116 ,
         \prgm_register/n1115 , \prgm_register/n1114 , \prgm_register/n1113 ,
         \prgm_register/n1112 , \prgm_register/n1111 , \prgm_register/n1110 ,
         \prgm_register/n1109 , \prgm_register/n1108 , \prgm_register/n1107 ,
         \prgm_register/n1106 , \prgm_register/n1105 , \prgm_register/n1104 ,
         \prgm_register/n1103 , \prgm_register/n1102 , \prgm_register/n1101 ,
         \prgm_register/n1100 , \prgm_register/n1099 , \prgm_register/n1098 ,
         \prgm_register/n1097 , \prgm_register/n1096 , \prgm_register/n1095 ,
         \prgm_register/n1094 , \prgm_register/n1093 , \prgm_register/n1092 ,
         \prgm_register/n1091 , \prgm_register/n1090 , \prgm_register/n1089 ,
         \prgm_register/n1088 , \prgm_register/n1087 , \prgm_register/n1086 ,
         \prgm_register/n1085 , \prgm_register/n1084 , \prgm_register/n1083 ,
         \prgm_register/n1082 , \prgm_register/n1081 , \prgm_register/n1080 ,
         \prgm_register/n1079 , \prgm_register/n1078 , \prgm_register/n1077 ,
         \prgm_register/n1076 , \prgm_register/n1075 , \prgm_register/n1074 ,
         \prgm_register/n1073 , \prgm_register/n1072 , \prgm_register/n1071 ,
         \prgm_register/n1070 , \prgm_register/n1069 , \prgm_register/n1068 ,
         \prgm_register/n1067 , \prgm_register/n1066 , \prgm_register/n1065 ,
         \prgm_register/n1064 , \prgm_register/n1063 , \prgm_register/n1062 ,
         \prgm_register/n1061 , \prgm_register/n1060 , \prgm_register/n1059 ,
         \prgm_register/n1058 , \prgm_register/n1057 , \prgm_register/n1056 ,
         \prgm_register/n1055 , \prgm_register/n1054 , \prgm_register/n1053 ,
         \prgm_register/n1052 , \prgm_register/n1051 , \prgm_register/n1050 ,
         \prgm_register/n1049 , \prgm_register/n1048 , \prgm_register/n1047 ,
         \prgm_register/n1046 , \prgm_register/n1045 , \prgm_register/n1044 ,
         \prgm_register/n1043 , \prgm_register/n1042 , \prgm_register/n1041 ,
         \prgm_register/n1040 , \prgm_register/n1039 , \prgm_register/n1038 ,
         \prgm_register/n1037 , \prgm_register/n1036 , \prgm_register/n1035 ,
         \prgm_register/n1034 , \prgm_register/n1033 , \prgm_register/n1032 ,
         \prgm_register/n1031 , \prgm_register/n1030 , \prgm_register/n1029 ,
         \prgm_register/n1028 , \prgm_register/n1027 , \prgm_register/n1026 ,
         \prgm_register/n1025 , \prgm_register/n1024 , \prgm_register/n1023 ,
         \prgm_register/n1022 , \prgm_register/n1021 , \prgm_register/n1020 ,
         \prgm_register/n1019 , \prgm_register/n1018 , \prgm_register/n1017 ,
         \prgm_register/n1016 , \prgm_register/n1015 , \prgm_register/n1014 ,
         \prgm_register/n1013 , \prgm_register/n1012 , \prgm_register/n1011 ,
         \prgm_register/n1010 , \prgm_register/n1009 , \prgm_register/n1008 ,
         \prgm_register/n1007 , \prgm_register/n1006 , \prgm_register/n1005 ,
         \prgm_register/n1004 , \prgm_register/n1003 , \prgm_register/n1002 ,
         \prgm_register/n1001 , \prgm_register/n1000 , \prgm_register/n999 ,
         \prgm_register/n998 , \prgm_register/n997 , \prgm_register/n996 ,
         \prgm_register/n995 , \prgm_register/n994 , \prgm_register/n993 ,
         \prgm_register/n992 , \prgm_register/n991 , \prgm_register/n990 ,
         \prgm_register/n989 , \prgm_register/n988 , \prgm_register/n987 ,
         \prgm_register/n986 , \prgm_register/n985 , \prgm_register/n984 ,
         \prgm_register/n983 , \prgm_register/n982 , \prgm_register/n981 ,
         \prgm_register/n980 , \prgm_register/n979 , \prgm_register/n978 ,
         \prgm_register/n977 , \prgm_register/n976 , \prgm_register/n975 ,
         \prgm_register/n974 , \prgm_register/n973 , \prgm_register/n972 ,
         \prgm_register/n971 , \prgm_register/n970 , \prgm_register/n969 ,
         \prgm_register/n968 , \prgm_register/n967 , \prgm_register/n966 ,
         \prgm_register/n965 , \prgm_register/n964 , \prgm_register/n963 ,
         \prgm_register/n962 , \prgm_register/n961 , \prgm_register/n960 ,
         \prgm_register/n959 , \prgm_register/n958 , \prgm_register/n957 ,
         \prgm_register/n956 , \prgm_register/n955 , \prgm_register/n954 ,
         \prgm_register/n953 , \prgm_register/n952 , \prgm_register/n951 ,
         \prgm_register/n950 , \prgm_register/n949 , \prgm_register/n948 ,
         \prgm_register/n947 , \prgm_register/n946 , \prgm_register/n945 ,
         \prgm_register/n944 , \prgm_register/n943 , \prgm_register/n942 ,
         \prgm_register/n941 , \prgm_register/n940 , \prgm_register/n939 ,
         \prgm_register/n938 , \prgm_register/n937 , \prgm_register/n936 ,
         \prgm_register/n935 , \prgm_register/n934 , \prgm_register/n933 ,
         \prgm_register/n932 , \prgm_register/n931 , \prgm_register/n930 ,
         \prgm_register/n929 , \prgm_register/n928 , \prgm_register/n927 ,
         \prgm_register/n926 , \prgm_register/n925 , \prgm_register/n924 ,
         \prgm_register/n923 , \prgm_register/n922 , \prgm_register/n921 ,
         \prgm_register/n920 , \prgm_register/n919 , \prgm_register/n918 ,
         \prgm_register/n917 , \prgm_register/n916 , \prgm_register/n915 ,
         \prgm_register/n914 , \prgm_register/n913 , \prgm_register/n912 ,
         \prgm_register/n911 , \prgm_register/n910 , \prgm_register/n909 ,
         \prgm_register/n908 , \prgm_register/n907 , \prgm_register/n906 ,
         \prgm_register/n905 , \prgm_register/n904 , \prgm_register/n903 ,
         \prgm_register/n902 , \prgm_register/n901 , \prgm_register/n900 ,
         \prgm_register/n899 , \prgm_register/n898 , \prgm_register/n897 ,
         \prgm_register/n896 , \prgm_register/n895 , \prgm_register/n894 ,
         \prgm_register/n893 , \prgm_register/n892 , \prgm_register/n891 ,
         \prgm_register/n890 , \prgm_register/n889 , \prgm_register/n888 ,
         \prgm_register/n887 , \prgm_register/n886 , \prgm_register/n885 ,
         \prgm_register/n884 , \prgm_register/n883 , \prgm_register/n882 ,
         \prgm_register/n881 , \prgm_register/n880 , \prgm_register/n879 ,
         \prgm_register/n878 , \prgm_register/n877 , \prgm_register/n876 ,
         \prgm_register/n875 , \prgm_register/n874 , \prgm_register/n873 ,
         \prgm_register/n872 , \prgm_register/n871 , \prgm_register/n870 ,
         \prgm_register/n869 , \prgm_register/n868 , \prgm_register/n867 ,
         \prgm_register/n866 , \prgm_register/n865 , \prgm_register/n864 ,
         \prgm_register/n863 , \prgm_register/n862 , \prgm_register/n861 ,
         \prgm_register/n860 , \prgm_register/n859 , \prgm_register/n858 ,
         \prgm_register/n857 , \prgm_register/n856 , \prgm_register/n855 ,
         \prgm_register/n854 , \prgm_register/n853 , \prgm_register/n852 ,
         \prgm_register/n851 , \prgm_register/n850 , \prgm_register/n849 ,
         \prgm_register/n848 , \prgm_register/n847 , \prgm_register/n846 ,
         \prgm_register/n845 , \prgm_register/n844 , \prgm_register/n843 ,
         \prgm_register/n842 , \prgm_register/n841 , \prgm_register/n840 ,
         \prgm_register/n839 , \prgm_register/n838 , \prgm_register/n837 ,
         \prgm_register/n836 , \prgm_register/n835 , \prgm_register/n834 ,
         \prgm_register/n833 , \prgm_register/n832 , \prgm_register/n831 ,
         \prgm_register/n830 , \prgm_register/n829 , \prgm_register/n828 ,
         \prgm_register/n827 , \prgm_register/n826 , \prgm_register/n825 ,
         \prgm_register/n824 , \prgm_register/n823 , \prgm_register/n822 ,
         \prgm_register/n821 , \prgm_register/n820 , \prgm_register/n819 ,
         \prgm_register/n818 , \prgm_register/n817 , \prgm_register/n816 ,
         \prgm_register/n815 , \prgm_register/n814 , \prgm_register/n813 ,
         \prgm_register/n812 , \prgm_register/n811 , \prgm_register/n810 ,
         \prgm_register/n809 , \prgm_register/n808 , \prgm_register/n807 ,
         \prgm_register/n806 , \prgm_register/n805 , \prgm_register/n804 ,
         \prgm_register/n803 , \prgm_register/n802 , \prgm_register/n801 ,
         \prgm_register/n800 , \prgm_register/n799 , \prgm_register/n798 ,
         \prgm_register/n797 , \prgm_register/n796 , \prgm_register/n795 ,
         \prgm_register/n794 , \prgm_register/n793 , \prgm_register/n792 ,
         \prgm_register/n791 , \prgm_register/n790 , \prgm_register/n789 ,
         \prgm_register/n788 , \prgm_register/n787 , \prgm_register/n786 ,
         \prgm_register/n785 , \prgm_register/n784 , \prgm_register/n783 ,
         \prgm_register/n782 , \prgm_register/n781 , \prgm_register/n780 ,
         \prgm_register/n779 , \prgm_register/n778 , \prgm_register/n777 ,
         \prgm_register/n776 , \prgm_register/n775 , \prgm_register/n774 ,
         \prgm_register/n773 , \prgm_register/n772 , \prgm_register/n771 ,
         \prgm_register/n770 , \prgm_register/n769 , \prgm_register/n768 ,
         \prgm_register/n767 , \prgm_register/n766 , \prgm_register/n765 ,
         \prgm_register/n764 , \prgm_register/n763 , \prgm_register/n762 ,
         \prgm_register/n761 , \prgm_register/n760 , \prgm_register/n759 ,
         \prgm_register/n758 , \prgm_register/n757 , \prgm_register/n756 ,
         \prgm_register/n755 , \prgm_register/n754 , \prgm_register/n753 ,
         \prgm_register/n752 , \prgm_register/n751 , \prgm_register/n750 ,
         \prgm_register/n749 , \prgm_register/n748 , \prgm_register/n747 ,
         \prgm_register/n746 , \prgm_register/n745 , \prgm_register/n744 ,
         \prgm_register/n743 , \prgm_register/n742 , \prgm_register/n741 ,
         \prgm_register/n740 , \prgm_register/n739 , \prgm_register/n738 ,
         \prgm_register/n737 , \prgm_register/n736 , \prgm_register/n735 ,
         \prgm_register/n734 , \prgm_register/n733 , \prgm_register/n732 ,
         \prgm_register/n731 , \prgm_register/n730 , \prgm_register/n729 ,
         \prgm_register/n728 , \prgm_register/n727 , \prgm_register/n726 ,
         \prgm_register/n725 , \prgm_register/n724 , \prgm_register/n723 ,
         \prgm_register/n722 , \prgm_register/n721 , \prgm_register/n720 ,
         \prgm_register/n719 , \prgm_register/n718 , \prgm_register/n717 ,
         \prgm_register/n716 , \prgm_register/n715 , \prgm_register/n714 ,
         \prgm_register/n713 , \prgm_register/n712 , \prgm_register/n711 ,
         \prgm_register/n710 , \prgm_register/n709 , \prgm_register/n708 ,
         \prgm_register/n707 , \prgm_register/n706 , \prgm_register/n705 ,
         \prgm_register/n704 , \prgm_register/n703 , \prgm_register/n702 ,
         \prgm_register/n701 , \prgm_register/n700 , \prgm_register/n699 ,
         \prgm_register/n698 , \prgm_register/n697 , \prgm_register/n696 ,
         \prgm_register/n695 , \prgm_register/n694 , \prgm_register/n693 ,
         \prgm_register/n692 , \prgm_register/n691 , \prgm_register/n690 ,
         \prgm_register/n689 , \prgm_register/n688 , \prgm_register/n687 ,
         \prgm_register/n686 , \prgm_register/n685 , \prgm_register/n684 ,
         \prgm_register/n683 , \prgm_register/n682 , \prgm_register/n681 ,
         \prgm_register/n680 , \prgm_register/n679 , \prgm_register/n678 ,
         \prgm_register/n677 , \prgm_register/n676 , \prgm_register/n675 ,
         \prgm_register/n674 , \prgm_register/n673 , \prgm_register/n672 ,
         \prgm_register/n671 , \prgm_register/n670 , \prgm_register/n669 ,
         \prgm_register/n668 , \prgm_register/n667 , \prgm_register/n666 ,
         \prgm_register/n665 , \prgm_register/n664 , \prgm_register/n663 ,
         \prgm_register/n662 , \prgm_register/n661 , \prgm_register/n660 ,
         \prgm_register/n659 , \prgm_register/n658 , \prgm_register/n657 ,
         \prgm_register/n656 , \prgm_register/n655 , \prgm_register/n654 ,
         \prgm_register/n653 , \prgm_register/n652 , \prgm_register/n651 ,
         \prgm_register/n650 , \prgm_register/n649 , \prgm_register/n648 ,
         \prgm_register/n647 , \prgm_register/n646 , \prgm_register/n645 ,
         \prgm_register/n644 , \prgm_register/n643 , \prgm_register/n642 ,
         \prgm_register/n641 , \prgm_register/n640 , \prgm_register/n639 ,
         \prgm_register/n638 , \prgm_register/n637 , \prgm_register/n636 ,
         \prgm_register/n635 , \prgm_register/n634 , \prgm_register/n633 ,
         \prgm_register/n632 , \prgm_register/n631 , \prgm_register/n630 ,
         \prgm_register/n629 , \prgm_register/n628 , \prgm_register/n627 ,
         \prgm_register/n626 , \prgm_register/n625 , \prgm_register/n624 ,
         \prgm_register/n623 , \prgm_register/n622 , \prgm_register/n621 ,
         \prgm_register/n620 , \prgm_register/n619 , \prgm_register/n618 ,
         \prgm_register/n617 , \prgm_register/n616 , \prgm_register/n615 ,
         \prgm_register/n614 , \prgm_register/n613 , \prgm_register/n612 ,
         \prgm_register/n611 , \prgm_register/n610 , \prgm_register/n609 ,
         \prgm_register/n608 , \prgm_register/n607 , \prgm_register/n606 ,
         \prgm_register/n605 , \prgm_register/n604 , \prgm_register/n603 ,
         \prgm_register/n602 , \prgm_register/n601 , \prgm_register/n600 ,
         \prgm_register/n599 , \prgm_register/n598 , \prgm_register/n597 ,
         \prgm_register/n596 , \prgm_register/n595 , \prgm_register/n594 ,
         \prgm_register/n593 , \prgm_register/n592 , \prgm_register/n591 ,
         \prgm_register/n590 , \prgm_register/n589 , \prgm_register/n588 ,
         \prgm_register/n587 , \prgm_register/n586 , \prgm_register/n585 ,
         \prgm_register/n584 , \prgm_register/n583 , \prgm_register/n582 ,
         \prgm_register/n581 , \prgm_register/n580 , \prgm_register/n579 ,
         \prgm_register/n578 , \prgm_register/n577 , \prgm_register/n576 ,
         \prgm_register/n575 , \prgm_register/n574 , \prgm_register/n573 ,
         \prgm_register/n572 , \prgm_register/n571 , \prgm_register/n570 ,
         \prgm_register/n569 , \prgm_register/n568 , \prgm_register/n567 ,
         \prgm_register/n566 , \prgm_register/n565 , \prgm_register/n564 ,
         \prgm_register/n563 , \prgm_register/n562 , \prgm_register/n561 ,
         \prgm_register/n560 , \prgm_register/n559 , \prgm_register/n558 ,
         \prgm_register/n557 , \prgm_register/n556 , \prgm_register/n555 ,
         \prgm_register/n554 , \prgm_register/n553 , \prgm_register/n552 ,
         \prgm_register/n551 , \prgm_register/n550 , \prgm_register/n549 ,
         \prgm_register/n548 , \prgm_register/n547 , \prgm_register/n546 ,
         \prgm_register/n545 , \prgm_register/n544 , \prgm_register/n543 ,
         \prgm_register/n542 , \prgm_register/n541 , \prgm_register/n540 ,
         \prgm_register/n539 , \prgm_register/n538 , \prgm_register/n537 ,
         \prgm_register/n536 , \prgm_register/n535 , \prgm_register/n534 ,
         \prgm_register/n533 , \prgm_register/n532 , \prgm_register/n531 ,
         \prgm_register/n530 , \prgm_register/n529 , \prgm_register/n528 ,
         \prgm_register/n527 , \prgm_register/n526 , \prgm_register/n525 ,
         \prgm_register/n524 , \prgm_register/n523 , \prgm_register/n522 ,
         \prgm_register/n521 , \prgm_register/n520 , \prgm_register/n519 ,
         \prgm_register/n518 , \prgm_register/n517 , \prgm_register/n516 ,
         \prgm_register/n515 , \prgm_register/n514 , \prgm_register/n513 ,
         \prgm_register/n512 , \prgm_register/n511 , \prgm_register/n510 ,
         \prgm_register/n509 , \prgm_register/n508 , \prgm_register/n507 ,
         \prgm_register/n506 , \prgm_register/n505 , \prgm_register/n504 ,
         \prgm_register/n503 , \prgm_register/n502 , \prgm_register/n501 ,
         \prgm_register/n500 , \prgm_register/n499 , \prgm_register/n498 ,
         \prgm_register/n497 , \prgm_register/n496 , \prgm_register/n495 ,
         \prgm_register/n494 , \prgm_register/n493 , \prgm_register/n492 ,
         \prgm_register/n491 , \prgm_register/n490 , \prgm_register/n489 ,
         \prgm_register/n488 , \prgm_register/n487 , \prgm_register/n486 ,
         \prgm_register/n485 , \prgm_register/n484 , \prgm_register/n483 ,
         \prgm_register/n482 , \prgm_register/n481 , \prgm_register/n480 ,
         \prgm_register/n479 , \prgm_register/n478 , \prgm_register/n477 ,
         \prgm_register/n476 , \prgm_register/n475 , \prgm_register/n474 ,
         \prgm_register/n473 , \prgm_register/n472 , \prgm_register/n471 ,
         \prgm_register/n470 , \prgm_register/n469 , \prgm_register/n468 ,
         \prgm_register/n467 , \prgm_register/n466 , \prgm_register/n465 ,
         \prgm_register/n464 , \prgm_register/n463 , \prgm_register/n462 ,
         \prgm_register/n461 , \prgm_register/n460 , \prgm_register/n459 ,
         \prgm_register/n458 , \prgm_register/n457 , \prgm_register/n456 ,
         \prgm_register/n455 , \prgm_register/n454 , \prgm_register/n453 ,
         \prgm_register/n452 , \prgm_register/n451 , \prgm_register/n450 ,
         \prgm_register/n449 , \prgm_register/n448 , \prgm_register/n447 ,
         \prgm_register/n446 , \prgm_register/n445 , \prgm_register/n444 ,
         \prgm_register/n443 , \prgm_register/n442 , \prgm_register/n441 ,
         \prgm_register/n440 , \prgm_register/n439 , \prgm_register/n438 ,
         \prgm_register/n437 , \prgm_register/n436 , \prgm_register/n435 ,
         \prgm_register/n434 , \prgm_register/n433 , \prgm_register/n432 ,
         \prgm_register/n431 , \prgm_register/n430 , \prgm_register/n429 ,
         \prgm_register/n428 , \prgm_register/n427 , \prgm_register/n426 ,
         \prgm_register/n425 , \prgm_register/n424 , \prgm_register/n423 ,
         \prgm_register/n422 , \prgm_register/n421 , \prgm_register/n420 ,
         \prgm_register/n419 , \prgm_register/n418 , \prgm_register/n417 ,
         \prgm_register/n416 , \prgm_register/n415 , \prgm_register/n414 ,
         \prgm_register/n413 , \prgm_register/n412 , \prgm_register/n411 ,
         \prgm_register/n410 , \prgm_register/n409 , \prgm_register/n408 ,
         \prgm_register/n407 , \prgm_register/n406 , \prgm_register/n405 ,
         \prgm_register/n404 , \prgm_register/n403 , \prgm_register/n402 ,
         \prgm_register/n401 , \prgm_register/n400 , \prgm_register/n399 ,
         \prgm_register/n398 , \prgm_register/n397 , \prgm_register/n396 ,
         \prgm_register/n395 , \prgm_register/n394 , \prgm_register/n393 ,
         \prgm_register/n392 , \prgm_register/n391 , \prgm_register/n390 ,
         \prgm_register/n389 , \prgm_register/n388 , \prgm_register/n387 ,
         \prgm_register/n386 , \prgm_register/n385 , \prgm_register/n384 ,
         \prgm_register/n383 , \prgm_register/n382 , \prgm_register/n381 ,
         \prgm_register/n380 , \prgm_register/n379 , \prgm_register/n378 ,
         \prgm_register/n377 , \prgm_register/n376 , \prgm_register/n375 ,
         \prgm_register/n374 , \prgm_register/n373 , \prgm_register/n372 ,
         \prgm_register/n371 , \prgm_register/n370 , \prgm_register/n369 ,
         \prgm_register/n368 , \prgm_register/n367 , \prgm_register/n366 ,
         \prgm_register/n365 , \prgm_register/n364 , \prgm_register/n363 ,
         \prgm_register/n362 , \prgm_register/n361 , \prgm_register/n360 ,
         \prgm_register/n359 , \prgm_register/n358 , \prgm_register/n357 ,
         \prgm_register/n356 , \prgm_register/n355 , \prgm_register/n354 ,
         \prgm_register/n353 , \prgm_register/n352 , \prgm_register/n351 ,
         \prgm_register/n350 , \prgm_register/n349 , \prgm_register/n348 ,
         \prgm_register/n347 , \prgm_register/n346 , \prgm_register/n345 ,
         \prgm_register/n344 , \prgm_register/n343 , \prgm_register/n342 ,
         \prgm_register/n341 , \prgm_register/n340 , \prgm_register/n339 ,
         \prgm_register/n338 , \prgm_register/n337 , \prgm_register/n336 ,
         \prgm_register/n335 , \prgm_register/n334 , \prgm_register/n333 ,
         \prgm_register/n332 , \prgm_register/n331 , \prgm_register/n330 ,
         \prgm_register/n329 , \prgm_register/n328 , \prgm_register/n327 ,
         \prgm_register/n326 , \prgm_register/n325 , \prgm_register/n324 ,
         \prgm_register/n323 , \prgm_register/n322 , \prgm_register/n321 ,
         \prgm_register/n320 , \prgm_register/n319 , \prgm_register/n318 ,
         \prgm_register/n317 , \prgm_register/n316 , \prgm_register/n315 ,
         \prgm_register/n314 , \prgm_register/n313 , \prgm_register/n312 ,
         \prgm_register/n311 , \prgm_register/n310 , \prgm_register/n309 ,
         \prgm_register/n308 , \prgm_register/n307 , \prgm_register/n306 ,
         \prgm_register/n305 , \prgm_register/n304 , \prgm_register/n303 ,
         \prgm_register/n302 , \prgm_register/n301 , \prgm_register/n300 ,
         \prgm_register/n299 , \prgm_register/n298 , \prgm_register/n297 ,
         \prgm_register/n296 , \prgm_register/n295 , \prgm_register/n294 ,
         \prgm_register/n293 , \prgm_register/n292 , \prgm_register/n291 ,
         \prgm_register/n290 , \prgm_register/n289 , \prgm_register/n288 ,
         \prgm_register/n287 , \prgm_register/n286 , \prgm_register/n285 ,
         \prgm_register/n284 , \prgm_register/n283 , \prgm_register/n282 ,
         \prgm_register/n281 , \prgm_register/n280 , \prgm_register/n279 ,
         \prgm_register/n278 , \prgm_register/n277 , \prgm_register/n276 ,
         \prgm_register/n275 , \prgm_register/n274 , \prgm_register/n273 ,
         \prgm_register/n272 , \prgm_register/n271 , \prgm_register/n270 ,
         \prgm_register/n269 , \prgm_register/n268 , \prgm_register/n267 ,
         \prgm_register/n266 , \prgm_register/n265 , \prgm_register/n264 ,
         \prgm_register/n263 , \prgm_register/n262 , \prgm_register/n261 ,
         \prgm_register/n260 , \prgm_register/n259 , \prgm_register/n258 ,
         \prgm_register/n257 , \prgm_register/n256 , \prgm_register/n255 ,
         \prgm_register/n254 , \prgm_register/n253 , \prgm_register/n252 ,
         \prgm_register/n251 , \prgm_register/n250 , \prgm_register/n249 ,
         \prgm_register/n248 , \prgm_register/n247 , \prgm_register/n246 ,
         \prgm_register/n245 , \prgm_register/n244 , \prgm_register/n243 ,
         \prgm_register/n242 , \prgm_register/n241 , \prgm_register/n240 ,
         \prgm_register/n239 , \prgm_register/n238 , \prgm_register/n237 ,
         \prgm_register/n236 , \prgm_register/n235 , \prgm_register/n234 ,
         \prgm_register/n233 , \prgm_register/n232 , \prgm_register/n231 ,
         \prgm_register/n230 , \prgm_register/n229 , \prgm_register/n228 ,
         \prgm_register/n227 , \prgm_register/n226 , \prgm_register/n225 ,
         \prgm_register/n224 , \prgm_register/n223 , \prgm_register/n222 ,
         \prgm_register/n221 , \prgm_register/n220 , \prgm_register/n219 ,
         \prgm_register/n218 , \prgm_register/n217 , \prgm_register/n216 ,
         \prgm_register/n215 , \prgm_register/n214 , \prgm_register/n213 ,
         \prgm_register/n212 , \prgm_register/n211 , \prgm_register/n210 ,
         \prgm_register/n209 , \prgm_register/n208 , \prgm_register/n207 ,
         \prgm_register/n206 , \prgm_register/n205 , \prgm_register/n204 ,
         \prgm_register/n203 , \prgm_register/n202 , \prgm_register/n201 ,
         \prgm_register/n200 , \prgm_register/n199 , \prgm_register/n198 ,
         \prgm_register/n197 , \prgm_register/n196 , \prgm_register/n195 ,
         \prgm_register/n194 , \prgm_register/n193 , \prgm_register/n192 ,
         \prgm_register/n191 , \prgm_register/n190 , \prgm_register/n189 ,
         \prgm_register/n188 , \prgm_register/n187 , \prgm_register/n186 ,
         \prgm_register/n185 , \prgm_register/n184 , \prgm_register/n183 ,
         \prgm_register/n182 , \prgm_register/n181 , \prgm_register/n180 ,
         \prgm_register/n179 , \prgm_register/n178 , \prgm_register/n177 ,
         \prgm_register/n176 , \prgm_register/n175 , \prgm_register/n174 ,
         \prgm_register/n173 , \prgm_register/n172 , \prgm_register/n171 ,
         \prgm_register/n170 , \prgm_register/n169 , \prgm_register/n168 ,
         \prgm_register/n167 , \prgm_register/n166 , \prgm_register/n165 ,
         \prgm_register/n164 , \prgm_register/n163 , \prgm_register/n162 ,
         \prgm_register/n161 , \prgm_register/n160 , \prgm_register/n159 ,
         \prgm_register/n158 , \prgm_register/n157 , \prgm_register/n156 ,
         \prgm_register/n155 , \prgm_register/n154 , \prgm_register/n153 ,
         \prgm_register/n152 , \prgm_register/n151 , \prgm_register/n150 ,
         \prgm_register/n149 , \prgm_register/n148 , \prgm_register/n147 ,
         \prgm_register/n146 , \prgm_register/n145 , \prgm_register/n144 ,
         \prgm_register/n143 , \prgm_register/n142 , \prgm_register/n141 ,
         \prgm_register/n140 , \prgm_register/n139 , \prgm_register/n138 ,
         \prgm_register/n137 , \prgm_register/n136 , \prgm_register/n135 ,
         \prgm_register/n134 , \prgm_register/n133 , \prgm_register/n132 ,
         \prgm_register/n131 , \prgm_register/n130 , \prgm_register/n129 ,
         \prgm_register/n128 , \prgm_register/n127 , \prgm_register/n126 ,
         \prgm_register/n125 , \prgm_register/n124 , \prgm_register/n123 ,
         \prgm_register/n122 , \prgm_register/n121 , \prgm_register/n120 ,
         \prgm_register/n119 , \prgm_register/n118 , \prgm_register/n117 ,
         \prgm_register/n116 , \prgm_register/n115 , \prgm_register/n114 ,
         \prgm_register/n113 , \prgm_register/n112 , \prgm_register/n111 ,
         \prgm_register/n110 , \prgm_register/n109 , \prgm_register/n108 ,
         \prgm_register/n107 , \prgm_register/n106 , \prgm_register/n105 ,
         \prgm_register/n104 , \prgm_register/n103 , \prgm_register/n102 ,
         \prgm_register/n101 , \prgm_register/n100 , \prgm_register/n99 ,
         \prgm_register/n98 , \prgm_register/n97 , \prgm_register/n96 ,
         \prgm_register/n95 , \prgm_register/n94 , \prgm_register/n93 ,
         \prgm_register/n92 , \prgm_register/n91 , \prgm_register/n90 ,
         \prgm_register/n89 , \prgm_register/n88 , \prgm_register/n87 ,
         \prgm_register/n86 , \prgm_register/n85 , \prgm_register/n84 ,
         \prgm_register/n83 , \prgm_register/n82 , \prgm_register/n81 ,
         \prgm_register/n80 , \prgm_register/n79 , \prgm_register/n78 ,
         \prgm_register/n77 , \prgm_register/n76 , \prgm_register/n75 ,
         \prgm_register/n74 , \prgm_register/n73 , \prgm_register/n72 ,
         \prgm_register/n71 , \prgm_register/n70 , \prgm_register/n69 ,
         \prgm_register/n68 , \prgm_register/n67 , \prgm_register/n66 ,
         \prgm_register/n65 , \prgm_register/n64 , \prgm_register/n63 ,
         \prgm_register/n62 , \prgm_register/n61 , \prgm_register/n60 ,
         \prgm_register/n59 , \prgm_register/n58 , \prgm_register/n57 ,
         \prgm_register/n56 , \prgm_register/n55 , \prgm_register/n54 ,
         \prgm_register/n53 , \prgm_register/n52 , \prgm_register/n51 ,
         \prgm_register/n50 , \prgm_register/n49 , \prgm_register/n48 ,
         \prgm_register/n47 , \prgm_register/n46 , \prgm_register/n45 ,
         \prgm_register/n44 , \prgm_register/n43 , \prgm_register/n42 ,
         \prgm_register/n41 , \prgm_register/n40 , \prgm_register/n39 ,
         \prgm_register/n38 , \prgm_register/n37 , \prgm_register/n36 ,
         \prgm_register/n35 , \prgm_register/n34 , \prgm_register/n33 ,
         \prgm_register/n32 , \prgm_register/n31 , \prgm_register/n30 ,
         \prgm_register/n29 , \prgm_register/n28 , \prgm_register/n27 ,
         \prgm_register/n26 , \prgm_register/n25 , \prgm_register/n24 ,
         \prgm_register/n23 , \prgm_register/n22 , \prgm_register/n21 ,
         \prgm_register/n20 , \prgm_register/n19 , \prgm_register/n18 ,
         \prgm_register/n17 , \prgm_register/n16 , \prgm_register/n15 ,
         \prgm_register/n14 , \prgm_register/n13 , \prgm_register/n12 ,
         \prgm_register/n11 , \prgm_register/n10 , \prgm_register/n9 ,
         \prgm_register/n8 , \prgm_register/n7 , \prgm_register/n6 ,
         \prgm_register/n5 , \prgm_register/n4 , \prgm_register/n3 ,
         \prgm_register/n2 , \prgm_register/n1 , \prgm_register/en_not ,
         \prgm_register/clear_not , \comparator/n2046 , \comparator/n2045 ,
         \comparator/n2044 , \comparator/n2043 , \comparator/n2042 ,
         \comparator/n2041 , \comparator/n2040 , \comparator/n2039 ,
         \comparator/n2038 , \comparator/n2037 , \comparator/n2036 ,
         \comparator/n2035 , \comparator/n2034 , \comparator/n2033 ,
         \comparator/n2032 , \comparator/n2031 , \comparator/n2030 ,
         \comparator/n2029 , \comparator/n2028 , \comparator/n2027 ,
         \comparator/n2026 , \comparator/n2025 , \comparator/n2024 ,
         \comparator/n2023 , \comparator/n2022 , \comparator/n2021 ,
         \comparator/n2020 , \comparator/n2019 , \comparator/n2018 ,
         \comparator/n2017 , \comparator/n2016 , \comparator/n2015 ,
         \comparator/n2014 , \comparator/n2013 , \comparator/n2012 ,
         \comparator/n2011 , \comparator/n2010 , \comparator/n2009 ,
         \comparator/n2008 , \comparator/n2007 , \comparator/n2006 ,
         \comparator/n2005 , \comparator/n2004 , \comparator/n2003 ,
         \comparator/n2002 , \comparator/n2001 , \comparator/n2000 ,
         \comparator/n1999 , \comparator/n1998 , \comparator/n1997 ,
         \comparator/n1996 , \comparator/n1995 , \comparator/n1994 ,
         \comparator/n1993 , \comparator/n1992 , \comparator/n1991 ,
         \comparator/n1990 , \comparator/n1989 , \comparator/n1988 ,
         \comparator/n1987 , \comparator/n1986 , \comparator/n1985 ,
         \comparator/n1984 , \comparator/n1983 , \comparator/n1982 ,
         \comparator/n1981 , \comparator/n1980 , \comparator/n1979 ,
         \comparator/n1978 , \comparator/n1977 , \comparator/n1976 ,
         \comparator/n1975 , \comparator/n1974 , \comparator/n1973 ,
         \comparator/n1972 , \comparator/n1971 , \comparator/n1970 ,
         \comparator/n1969 , \comparator/n1968 , \comparator/n1967 ,
         \comparator/n1966 , \comparator/n1965 , \comparator/n1964 ,
         \comparator/n1963 , \comparator/n1962 , \comparator/n1961 ,
         \comparator/n1960 , \comparator/n1959 , \comparator/n1958 ,
         \comparator/n1957 , \comparator/n1956 , \comparator/n1955 ,
         \comparator/n1954 , \comparator/n1953 , \comparator/n1952 ,
         \comparator/n1951 , \comparator/n1950 , \comparator/n1949 ,
         \comparator/n1948 , \comparator/n1947 , \comparator/n1946 ,
         \comparator/n1945 , \comparator/n1944 , \comparator/n1943 ,
         \comparator/n1942 , \comparator/n1941 , \comparator/n1940 ,
         \comparator/n1939 , \comparator/n1938 , \comparator/n1937 ,
         \comparator/n1936 , \comparator/n1935 , \comparator/n1934 ,
         \comparator/n1933 , \comparator/n1932 , \comparator/n1931 ,
         \comparator/n1930 , \comparator/n1929 , \comparator/n1928 ,
         \comparator/n1927 , \comparator/n1926 , \comparator/n1925 ,
         \comparator/n1924 , \comparator/n1923 , \comparator/n1922 ,
         \comparator/n1921 , \comparator/n1920 , \comparator/n1919 ,
         \comparator/n1918 , \comparator/n1917 , \comparator/n1916 ,
         \comparator/n1915 , \comparator/n1914 , \comparator/n1913 ,
         \comparator/n1912 , \comparator/n1911 , \comparator/n1910 ,
         \comparator/n1909 , \comparator/n1908 , \comparator/n1907 ,
         \comparator/n1906 , \comparator/n1905 , \comparator/n1904 ,
         \comparator/n1903 , \comparator/n1902 , \comparator/n1901 ,
         \comparator/n1900 , \comparator/n1899 , \comparator/n1898 ,
         \comparator/n1897 , \comparator/n1896 , \comparator/n1895 ,
         \comparator/n1894 , \comparator/n1893 , \comparator/n1892 ,
         \comparator/n1891 , \comparator/n1890 , \comparator/n1889 ,
         \comparator/n1888 , \comparator/n1887 , \comparator/n1886 ,
         \comparator/n1885 , \comparator/n1884 , \comparator/n1883 ,
         \comparator/n1882 , \comparator/n1881 , \comparator/n1880 ,
         \comparator/n1879 , \comparator/n1878 , \comparator/n1877 ,
         \comparator/n1876 , \comparator/n1875 , \comparator/n1874 ,
         \comparator/n1873 , \comparator/n1872 , \comparator/n1871 ,
         \comparator/n1870 , \comparator/n1869 , \comparator/n1868 ,
         \comparator/n1867 , \comparator/n1866 , \comparator/n1865 ,
         \comparator/n1864 , \comparator/n1863 , \comparator/n1862 ,
         \comparator/n1861 , \comparator/n1860 , \comparator/n1859 ,
         \comparator/n1858 , \comparator/n1857 , \comparator/n1856 ,
         \comparator/n1855 , \comparator/n1854 , \comparator/n1853 ,
         \comparator/n1852 , \comparator/n1851 , \comparator/n1850 ,
         \comparator/n1849 , \comparator/n1848 , \comparator/n1847 ,
         \comparator/n1846 , \comparator/n1845 , \comparator/n1844 ,
         \comparator/n1843 , \comparator/n1842 , \comparator/n1841 ,
         \comparator/n1840 , \comparator/n1839 , \comparator/n1838 ,
         \comparator/n1837 , \comparator/n1836 , \comparator/n1835 ,
         \comparator/n1834 , \comparator/n1833 , \comparator/n1832 ,
         \comparator/n1831 , \comparator/n1830 , \comparator/n1829 ,
         \comparator/n1828 , \comparator/n1827 , \comparator/n1826 ,
         \comparator/n1825 , \comparator/n1824 , \comparator/n1823 ,
         \comparator/n1822 , \comparator/n1821 , \comparator/n1820 ,
         \comparator/n1819 , \comparator/n1818 , \comparator/n1817 ,
         \comparator/n1816 , \comparator/n1815 , \comparator/n1814 ,
         \comparator/n1813 , \comparator/n1812 , \comparator/n1811 ,
         \comparator/n1810 , \comparator/n1809 , \comparator/n1808 ,
         \comparator/n1807 , \comparator/n1806 , \comparator/n1805 ,
         \comparator/n1804 , \comparator/n1803 , \comparator/n1802 ,
         \comparator/n1801 , \comparator/n1800 , \comparator/n1799 ,
         \comparator/n1798 , \comparator/n1797 , \comparator/n1796 ,
         \comparator/n1795 , \comparator/n1794 , \comparator/n1793 ,
         \comparator/n1792 , \comparator/n1791 , \comparator/n1790 ,
         \comparator/n1789 , \comparator/n1788 , \comparator/n1787 ,
         \comparator/n1786 , \comparator/n1785 , \comparator/n1784 ,
         \comparator/n1783 , \comparator/n1782 , \comparator/n1781 ,
         \comparator/n1780 , \comparator/n1779 , \comparator/n1778 ,
         \comparator/n1777 , \comparator/n1776 , \comparator/n1775 ,
         \comparator/n1774 , \comparator/n1773 , \comparator/n1772 ,
         \comparator/n1771 , \comparator/n1770 , \comparator/n1769 ,
         \comparator/n1768 , \comparator/n1767 , \comparator/n1766 ,
         \comparator/n1765 , \comparator/n1764 , \comparator/n1763 ,
         \comparator/n1762 , \comparator/n1761 , \comparator/n1760 ,
         \comparator/n1759 , \comparator/n1758 , \comparator/n1757 ,
         \comparator/n1756 , \comparator/n1755 , \comparator/n1754 ,
         \comparator/n1753 , \comparator/n1752 , \comparator/n1751 ,
         \comparator/n1750 , \comparator/n1749 , \comparator/n1748 ,
         \comparator/n1747 , \comparator/n1746 , \comparator/n1745 ,
         \comparator/n1744 , \comparator/n1743 , \comparator/n1742 ,
         \comparator/n1741 , \comparator/n1740 , \comparator/n1739 ,
         \comparator/n1738 , \comparator/n1737 , \comparator/n1736 ,
         \comparator/n1735 , \comparator/n1734 , \comparator/n1733 ,
         \comparator/n1732 , \comparator/n1731 , \comparator/n1730 ,
         \comparator/n1729 , \comparator/n1728 , \comparator/n1727 ,
         \comparator/n1726 , \comparator/n1725 , \comparator/n1724 ,
         \comparator/n1723 , \comparator/n1722 , \comparator/n1721 ,
         \comparator/n1720 , \comparator/n1719 , \comparator/n1718 ,
         \comparator/n1717 , \comparator/n1716 , \comparator/n1715 ,
         \comparator/n1714 , \comparator/n1713 , \comparator/n1712 ,
         \comparator/n1711 , \comparator/n1710 , \comparator/n1709 ,
         \comparator/n1708 , \comparator/n1707 , \comparator/n1706 ,
         \comparator/n1705 , \comparator/n1704 , \comparator/n1703 ,
         \comparator/n1702 , \comparator/n1701 , \comparator/n1700 ,
         \comparator/n1699 , \comparator/n1698 , \comparator/n1697 ,
         \comparator/n1696 , \comparator/n1695 , \comparator/n1694 ,
         \comparator/n1693 , \comparator/n1692 , \comparator/n1691 ,
         \comparator/n1690 , \comparator/n1689 , \comparator/n1688 ,
         \comparator/n1687 , \comparator/n1686 , \comparator/n1685 ,
         \comparator/n1684 , \comparator/n1683 , \comparator/n1682 ,
         \comparator/n1681 , \comparator/n1680 , \comparator/n1679 ,
         \comparator/n1678 , \comparator/n1677 , \comparator/n1676 ,
         \comparator/n1675 , \comparator/n1674 , \comparator/n1673 ,
         \comparator/n1672 , \comparator/n1671 , \comparator/n1670 ,
         \comparator/n1669 , \comparator/n1668 , \comparator/n1667 ,
         \comparator/n1666 , \comparator/n1665 , \comparator/n1664 ,
         \comparator/n1663 , \comparator/n1662 , \comparator/n1661 ,
         \comparator/n1660 , \comparator/n1659 , \comparator/n1658 ,
         \comparator/n1657 , \comparator/n1656 , \comparator/n1655 ,
         \comparator/n1654 , \comparator/n1653 , \comparator/n1652 ,
         \comparator/n1651 , \comparator/n1650 , \comparator/n1649 ,
         \comparator/n1648 , \comparator/n1647 , \comparator/n1646 ,
         \comparator/n1645 , \comparator/n1644 , \comparator/n1643 ,
         \comparator/n1642 , \comparator/n1641 , \comparator/n1640 ,
         \comparator/n1639 , \comparator/n1638 , \comparator/n1637 ,
         \comparator/n1636 , \comparator/n1635 , \comparator/n1634 ,
         \comparator/n1633 , \comparator/n1632 , \comparator/n1631 ,
         \comparator/n1630 , \comparator/n1629 , \comparator/n1628 ,
         \comparator/n1627 , \comparator/n1626 , \comparator/n1625 ,
         \comparator/n1624 , \comparator/n1623 , \comparator/n1622 ,
         \comparator/n1621 , \comparator/n1620 , \comparator/n1619 ,
         \comparator/n1618 , \comparator/n1617 , \comparator/n1616 ,
         \comparator/n1615 , \comparator/n1614 , \comparator/n1613 ,
         \comparator/n1612 , \comparator/n1611 , \comparator/n1610 ,
         \comparator/n1609 , \comparator/n1608 , \comparator/n1607 ,
         \comparator/n1606 , \comparator/n1605 , \comparator/n1604 ,
         \comparator/n1603 , \comparator/n1602 , \comparator/n1601 ,
         \comparator/n1600 , \comparator/n1599 , \comparator/n1598 ,
         \comparator/n1597 , \comparator/n1596 , \comparator/n1595 ,
         \comparator/n1594 , \comparator/n1593 , \comparator/n1592 ,
         \comparator/n1591 , \comparator/n1590 , \comparator/n1589 ,
         \comparator/n1588 , \comparator/n1587 , \comparator/n1586 ,
         \comparator/n1585 , \comparator/n1584 , \comparator/n1583 ,
         \comparator/n1582 , \comparator/n1581 , \comparator/n1580 ,
         \comparator/n1579 , \comparator/n1578 , \comparator/n1577 ,
         \comparator/n1576 , \comparator/n1575 , \comparator/n1574 ,
         \comparator/n1573 , \comparator/n1572 , \comparator/n1571 ,
         \comparator/n1570 , \comparator/n1569 , \comparator/n1568 ,
         \comparator/n1567 , \comparator/n1566 , \comparator/n1565 ,
         \comparator/n1564 , \comparator/n1563 , \comparator/n1562 ,
         \comparator/n1561 , \comparator/n1560 , \comparator/n1559 ,
         \comparator/n1558 , \comparator/n1557 , \comparator/n1556 ,
         \comparator/n1555 , \comparator/n1554 , \comparator/n1553 ,
         \comparator/n1552 , \comparator/n1551 , \comparator/n1550 ,
         \comparator/n1549 , \comparator/n1548 , \comparator/n1547 ,
         \comparator/n1546 , \comparator/n1545 , \comparator/n1544 ,
         \comparator/n1543 , \comparator/n1542 , \comparator/n1541 ,
         \comparator/n1540 , \comparator/n1539 , \comparator/n1538 ,
         \comparator/n1537 , \comparator/n1536 , \comparator/n1535 ,
         \comparator/n1534 , \comparator/n1533 , \comparator/n1532 ,
         \comparator/n1531 , \comparator/n1530 , \comparator/n1529 ,
         \comparator/n1528 , \comparator/n1527 , \comparator/n1526 ,
         \comparator/n1525 , \comparator/n1524 , \comparator/n1523 ,
         \comparator/n1522 , \comparator/n1521 , \comparator/n1520 ,
         \comparator/n1519 , \comparator/n1518 , \comparator/n1517 ,
         \comparator/n1516 , \comparator/n1515 , \comparator/n1514 ,
         \comparator/n1513 , \comparator/n1512 , \comparator/n1511 ,
         \comparator/n1510 , \comparator/n1509 , \comparator/n1508 ,
         \comparator/n1507 , \comparator/n1506 , \comparator/n1505 ,
         \comparator/n1504 , \comparator/n1503 , \comparator/n1502 ,
         \comparator/n1501 , \comparator/n1500 , \comparator/n1499 ,
         \comparator/n1498 , \comparator/n1497 , \comparator/n1496 ,
         \comparator/n1495 , \comparator/n1494 , \comparator/n1493 ,
         \comparator/n1492 , \comparator/n1491 , \comparator/n1490 ,
         \comparator/n1489 , \comparator/n1488 , \comparator/n1487 ,
         \comparator/n1486 , \comparator/n1485 , \comparator/n1484 ,
         \comparator/n1483 , \comparator/n1482 , \comparator/n1481 ,
         \comparator/n1480 , \comparator/n1479 , \comparator/n1478 ,
         \comparator/n1477 , \comparator/n1476 , \comparator/n1475 ,
         \comparator/n1474 , \comparator/n1473 , \comparator/n1472 ,
         \comparator/n1471 , \comparator/n1470 , \comparator/n1469 ,
         \comparator/n1468 , \comparator/n1467 , \comparator/n1466 ,
         \comparator/n1465 , \comparator/n1464 , \comparator/n1463 ,
         \comparator/n1462 , \comparator/n1461 , \comparator/n1460 ,
         \comparator/n1459 , \comparator/n1458 , \comparator/n1457 ,
         \comparator/n1456 , \comparator/n1455 , \comparator/n1454 ,
         \comparator/n1453 , \comparator/n1452 , \comparator/n1451 ,
         \comparator/n1450 , \comparator/n1449 , \comparator/n1448 ,
         \comparator/n1447 , \comparator/n1446 , \comparator/n1445 ,
         \comparator/n1444 , \comparator/n1443 , \comparator/n1442 ,
         \comparator/n1441 , \comparator/n1440 , \comparator/n1439 ,
         \comparator/n1438 , \comparator/n1437 , \comparator/n1436 ,
         \comparator/n1435 , \comparator/n1434 , \comparator/n1433 ,
         \comparator/n1432 , \comparator/n1431 , \comparator/n1430 ,
         \comparator/n1429 , \comparator/n1428 , \comparator/n1427 ,
         \comparator/n1426 , \comparator/n1425 , \comparator/n1424 ,
         \comparator/n1423 , \comparator/n1422 , \comparator/n1421 ,
         \comparator/n1420 , \comparator/n1419 , \comparator/n1418 ,
         \comparator/n1417 , \comparator/n1416 , \comparator/n1415 ,
         \comparator/n1414 , \comparator/n1413 , \comparator/n1412 ,
         \comparator/n1411 , \comparator/n1410 , \comparator/n1409 ,
         \comparator/n1408 , \comparator/n1407 , \comparator/n1406 ,
         \comparator/n1405 , \comparator/n1404 , \comparator/n1403 ,
         \comparator/n1402 , \comparator/n1401 , \comparator/n1400 ,
         \comparator/n1399 , \comparator/n1398 , \comparator/n1397 ,
         \comparator/n1396 , \comparator/n1395 , \comparator/n1394 ,
         \comparator/n1393 , \comparator/n1392 , \comparator/n1391 ,
         \comparator/n1390 , \comparator/n1389 , \comparator/n1388 ,
         \comparator/n1387 , \comparator/n1386 , \comparator/n1385 ,
         \comparator/n1384 , \comparator/n1383 , \comparator/n1382 ,
         \comparator/n1381 , \comparator/n1380 , \comparator/n1379 ,
         \comparator/n1378 , \comparator/n1377 , \comparator/n1376 ,
         \comparator/n1375 , \comparator/n1374 , \comparator/n1373 ,
         \comparator/n1372 , \comparator/n1371 , \comparator/n1370 ,
         \comparator/n1369 , \comparator/n1368 , \comparator/n1367 ,
         \comparator/n1366 , \comparator/n1365 , \comparator/n1364 ,
         \comparator/n1363 , \comparator/n1362 , \comparator/n1361 ,
         \comparator/n1360 , \comparator/n1359 , \comparator/n1358 ,
         \comparator/n1357 , \comparator/n1356 , \comparator/n1355 ,
         \comparator/n1354 , \comparator/n1353 , \comparator/n1352 ,
         \comparator/n1351 , \comparator/n1350 , \comparator/n1349 ,
         \comparator/n1348 , \comparator/n1347 , \comparator/n1346 ,
         \comparator/n1345 , \comparator/n1344 , \comparator/n1343 ,
         \comparator/n1342 , \comparator/n1341 , \comparator/n1340 ,
         \comparator/n1339 , \comparator/n1338 , \comparator/n1337 ,
         \comparator/n1336 , \comparator/n1335 , \comparator/n1334 ,
         \comparator/n1333 , \comparator/n1332 , \comparator/n1331 ,
         \comparator/n1330 , \comparator/n1329 , \comparator/n1328 ,
         \comparator/n1327 , \comparator/n1326 , \comparator/n1325 ,
         \comparator/n1324 , \comparator/n1323 , \comparator/n1322 ,
         \comparator/n1321 , \comparator/n1320 , \comparator/n1319 ,
         \comparator/n1318 , \comparator/n1317 , \comparator/n1316 ,
         \comparator/n1315 , \comparator/n1314 , \comparator/n1313 ,
         \comparator/n1312 , \comparator/n1311 , \comparator/n1310 ,
         \comparator/n1309 , \comparator/n1308 , \comparator/n1307 ,
         \comparator/n1306 , \comparator/n1305 , \comparator/n1304 ,
         \comparator/n1303 , \comparator/n1302 , \comparator/n1301 ,
         \comparator/n1300 , \comparator/n1299 , \comparator/n1298 ,
         \comparator/n1297 , \comparator/n1296 , \comparator/n1295 ,
         \comparator/n1294 , \comparator/n1293 , \comparator/n1292 ,
         \comparator/n1291 , \comparator/n1290 , \comparator/n1289 ,
         \comparator/n1288 , \comparator/n1287 , \comparator/n1286 ,
         \comparator/n1285 , \comparator/n1284 , \comparator/n1283 ,
         \comparator/n1282 , \comparator/n1281 , \comparator/n1280 ,
         \comparator/n1279 , \comparator/n1278 , \comparator/n1277 ,
         \comparator/n1276 , \comparator/n1275 , \comparator/n1274 ,
         \comparator/n1273 , \comparator/n1272 , \comparator/n1271 ,
         \comparator/n1270 , \comparator/n1269 , \comparator/n1268 ,
         \comparator/n1267 , \comparator/n1266 , \comparator/n1265 ,
         \comparator/n1264 , \comparator/n1263 , \comparator/n1262 ,
         \comparator/n1261 , \comparator/n1260 , \comparator/n1259 ,
         \comparator/n1258 , \comparator/n1257 , \comparator/n1256 ,
         \comparator/n1255 , \comparator/n1254 , \comparator/n1253 ,
         \comparator/n1252 , \comparator/n1251 , \comparator/n1250 ,
         \comparator/n1249 , \comparator/n1248 , \comparator/n1247 ,
         \comparator/n1246 , \comparator/n1245 , \comparator/n1244 ,
         \comparator/n1243 , \comparator/n1242 , \comparator/n1241 ,
         \comparator/n1240 , \comparator/n1239 , \comparator/n1238 ,
         \comparator/n1237 , \comparator/n1236 , \comparator/n1235 ,
         \comparator/n1234 , \comparator/n1233 , \comparator/n1232 ,
         \comparator/n1231 , \comparator/n1230 , \comparator/n1229 ,
         \comparator/n1228 , \comparator/n1227 , \comparator/n1226 ,
         \comparator/n1225 , \comparator/n1224 , \comparator/n1223 ,
         \comparator/n1222 , \comparator/n1221 , \comparator/n1220 ,
         \comparator/n1219 , \comparator/n1218 , \comparator/n1217 ,
         \comparator/n1216 , \comparator/n1215 , \comparator/n1214 ,
         \comparator/n1213 , \comparator/n1212 , \comparator/n1211 ,
         \comparator/n1210 , \comparator/n1209 , \comparator/n1208 ,
         \comparator/n1207 , \comparator/n1206 , \comparator/n1205 ,
         \comparator/n1204 , \comparator/n1203 , \comparator/n1202 ,
         \comparator/n1201 , \comparator/n1200 , \comparator/n1199 ,
         \comparator/n1198 , \comparator/n1197 , \comparator/n1196 ,
         \comparator/n1195 , \comparator/n1194 , \comparator/n1193 ,
         \comparator/n1192 , \comparator/n1191 , \comparator/n1190 ,
         \comparator/n1189 , \comparator/n1188 , \comparator/n1187 ,
         \comparator/n1186 , \comparator/n1185 , \comparator/n1184 ,
         \comparator/n1183 , \comparator/n1182 , \comparator/n1181 ,
         \comparator/n1180 , \comparator/n1179 , \comparator/n1178 ,
         \comparator/n1177 , \comparator/n1176 , \comparator/n1175 ,
         \comparator/n1174 , \comparator/n1173 , \comparator/n1172 ,
         \comparator/n1171 , \comparator/n1170 , \comparator/n1169 ,
         \comparator/n1168 , \comparator/n1167 , \comparator/n1166 ,
         \comparator/n1165 , \comparator/n1164 , \comparator/n1163 ,
         \comparator/n1162 , \comparator/n1161 , \comparator/n1160 ,
         \comparator/n1159 , \comparator/n1158 , \comparator/n1157 ,
         \comparator/n1156 , \comparator/n1155 , \comparator/n1154 ,
         \comparator/n1153 , \comparator/n1152 , \comparator/n1151 ,
         \comparator/n1150 , \comparator/n1149 , \comparator/n1148 ,
         \comparator/n1147 , \comparator/n1146 , \comparator/n1145 ,
         \comparator/n1144 , \comparator/n1143 , \comparator/n1142 ,
         \comparator/n1141 , \comparator/n1140 , \comparator/n1139 ,
         \comparator/n1138 , \comparator/n1137 , \comparator/n1136 ,
         \comparator/n1135 , \comparator/n1134 , \comparator/n1133 ,
         \comparator/n1132 , \comparator/n1131 , \comparator/n1130 ,
         \comparator/n1129 , \comparator/n1128 , \comparator/n1127 ,
         \comparator/n1126 , \comparator/n1125 , \comparator/n1124 ,
         \comparator/n1123 , \comparator/n1122 , \comparator/n1121 ,
         \comparator/n1120 , \comparator/n1119 , \comparator/n1118 ,
         \comparator/n1117 , \comparator/n1116 , \comparator/n1115 ,
         \comparator/n1114 , \comparator/n1113 , \comparator/n1112 ,
         \comparator/n1111 , \comparator/n1110 , \comparator/n1109 ,
         \comparator/n1108 , \comparator/n1107 , \comparator/n1106 ,
         \comparator/n1105 , \comparator/n1104 , \comparator/n1103 ,
         \comparator/n1102 , \comparator/n1101 , \comparator/n1100 ,
         \comparator/n1099 , \comparator/n1098 , \comparator/n1097 ,
         \comparator/n1096 , \comparator/n1095 , \comparator/n1094 ,
         \comparator/n1093 , \comparator/n1092 , \comparator/n1091 ,
         \comparator/n1090 , \comparator/n1089 , \comparator/n1088 ,
         \comparator/n1087 , \comparator/n1086 , \comparator/n1085 ,
         \comparator/n1084 , \comparator/n1083 , \comparator/n1082 ,
         \comparator/n1081 , \comparator/n1080 , \comparator/n1079 ,
         \comparator/n1078 , \comparator/n1077 , \comparator/n1076 ,
         \comparator/n1075 , \comparator/n1074 , \comparator/n1073 ,
         \comparator/n1072 , \comparator/n1071 , \comparator/n1070 ,
         \comparator/n1069 , \comparator/n1068 , \comparator/n1067 ,
         \comparator/n1066 , \comparator/n1065 , \comparator/n1064 ,
         \comparator/n1063 , \comparator/n1062 , \comparator/n1061 ,
         \comparator/n1060 , \comparator/n1059 , \comparator/n1058 ,
         \comparator/n1057 , \comparator/n1056 , \comparator/n1055 ,
         \comparator/n1054 , \comparator/n1053 , \comparator/n1052 ,
         \comparator/n1051 , \comparator/n1050 , \comparator/n1049 ,
         \comparator/n1048 , \comparator/n1047 , \comparator/n1046 ,
         \comparator/n1045 , \comparator/n1044 , \comparator/n1043 ,
         \comparator/n1042 , \comparator/n1041 , \comparator/n1040 ,
         \comparator/n1039 , \comparator/n1038 , \comparator/n1037 ,
         \comparator/n1036 , \comparator/n1035 , \comparator/n1034 ,
         \comparator/n1033 , \comparator/n1032 , \comparator/n1031 ,
         \comparator/n1030 , \comparator/n1029 , \comparator/n1028 ,
         \comparator/n1027 , \comparator/n1026 , \comparator/n1025 ,
         \comparator/n1024 , \comparator/n1023 , \comparator/n1022 ,
         \comparator/n1021 , \comparator/n1020 , \comparator/n1019 ,
         \comparator/n1018 , \comparator/n1017 , \comparator/n1016 ,
         \comparator/n1015 , \comparator/n1014 , \comparator/n1013 ,
         \comparator/n1012 , \comparator/n1011 , \comparator/n1010 ,
         \comparator/n1009 , \comparator/n1008 , \comparator/n1007 ,
         \comparator/n1006 , \comparator/n1005 , \comparator/n1004 ,
         \comparator/n1003 , \comparator/n1002 , \comparator/n1001 ,
         \comparator/n1000 , \comparator/n999 , \comparator/n998 ,
         \comparator/n997 , \comparator/n996 , \comparator/n995 ,
         \comparator/n994 , \comparator/n993 , \comparator/n992 ,
         \comparator/n991 , \comparator/n990 , \comparator/n989 ,
         \comparator/n988 , \comparator/n987 , \comparator/n986 ,
         \comparator/n985 , \comparator/n984 , \comparator/n983 ,
         \comparator/n982 , \comparator/n981 , \comparator/n980 ,
         \comparator/n979 , \comparator/n978 , \comparator/n977 ,
         \comparator/n976 , \comparator/n975 , \comparator/n974 ,
         \comparator/n973 , \comparator/n972 , \comparator/n971 ,
         \comparator/n970 , \comparator/n969 , \comparator/n968 ,
         \comparator/n967 , \comparator/n966 , \comparator/n965 ,
         \comparator/n964 , \comparator/n963 , \comparator/n962 ,
         \comparator/n961 , \comparator/n960 , \comparator/n959 ,
         \comparator/n958 , \comparator/n957 , \comparator/n956 ,
         \comparator/n955 , \comparator/n954 , \comparator/n953 ,
         \comparator/n952 , \comparator/n951 , \comparator/n950 ,
         \comparator/n949 , \comparator/n948 , \comparator/n947 ,
         \comparator/n946 , \comparator/n945 , \comparator/n944 ,
         \comparator/n943 , \comparator/n942 , \comparator/n941 ,
         \comparator/n940 , \comparator/n939 , \comparator/n938 ,
         \comparator/n937 , \comparator/n936 , \comparator/n935 ,
         \comparator/n934 , \comparator/n933 , \comparator/n932 ,
         \comparator/n931 , \comparator/n930 , \comparator/n929 ,
         \comparator/n928 , \comparator/n927 , \comparator/n926 ,
         \comparator/n925 , \comparator/n924 , \comparator/n923 ,
         \comparator/n922 , \comparator/n921 , \comparator/n920 ,
         \comparator/n919 , \comparator/n918 , \comparator/n917 ,
         \comparator/n916 , \comparator/n915 , \comparator/n914 ,
         \comparator/n913 , \comparator/n912 , \comparator/n911 ,
         \comparator/n910 , \comparator/n909 , \comparator/n908 ,
         \comparator/n907 , \comparator/n906 , \comparator/n905 ,
         \comparator/n904 , \comparator/n903 , \comparator/n902 ,
         \comparator/n901 , \comparator/n900 , \comparator/n899 ,
         \comparator/n898 , \comparator/n897 , \comparator/n896 ,
         \comparator/n895 , \comparator/n894 , \comparator/n893 ,
         \comparator/n892 , \comparator/n891 , \comparator/n890 ,
         \comparator/n889 , \comparator/n888 , \comparator/n887 ,
         \comparator/n886 , \comparator/n885 , \comparator/n884 ,
         \comparator/n883 , \comparator/n882 , \comparator/n881 ,
         \comparator/n880 , \comparator/n879 , \comparator/n878 ,
         \comparator/n877 , \comparator/n876 , \comparator/n875 ,
         \comparator/n874 , \comparator/n873 , \comparator/n872 ,
         \comparator/n871 , \comparator/n870 , \comparator/n869 ,
         \comparator/n868 , \comparator/n867 , \comparator/n866 ,
         \comparator/n865 , \comparator/n864 , \comparator/n863 ,
         \comparator/n862 , \comparator/n861 , \comparator/n860 ,
         \comparator/n859 , \comparator/n858 , \comparator/n857 ,
         \comparator/n856 , \comparator/n855 , \comparator/n854 ,
         \comparator/n853 , \comparator/n852 , \comparator/n851 ,
         \comparator/n850 , \comparator/n849 , \comparator/n848 ,
         \comparator/n847 , \comparator/n846 , \comparator/n845 ,
         \comparator/n844 , \comparator/n843 , \comparator/n842 ,
         \comparator/n841 , \comparator/n840 , \comparator/n839 ,
         \comparator/n838 , \comparator/n837 , \comparator/n836 ,
         \comparator/n835 , \comparator/n834 , \comparator/n833 ,
         \comparator/n832 , \comparator/n831 , \comparator/n830 ,
         \comparator/n829 , \comparator/n828 , \comparator/n827 ,
         \comparator/n826 , \comparator/n825 , \comparator/n824 ,
         \comparator/n823 , \comparator/n822 , \comparator/n821 ,
         \comparator/n820 , \comparator/n819 , \comparator/n818 ,
         \comparator/n817 , \comparator/n816 , \comparator/n815 ,
         \comparator/n814 , \comparator/n813 , \comparator/n812 ,
         \comparator/n811 , \comparator/n810 , \comparator/n809 ,
         \comparator/n808 , \comparator/n807 , \comparator/n806 ,
         \comparator/n805 , \comparator/n804 , \comparator/n803 ,
         \comparator/n802 , \comparator/n801 , \comparator/n800 ,
         \comparator/n799 , \comparator/n798 , \comparator/n797 ,
         \comparator/n796 , \comparator/n795 , \comparator/n794 ,
         \comparator/n793 , \comparator/n792 , \comparator/n791 ,
         \comparator/n790 , \comparator/n789 , \comparator/n788 ,
         \comparator/n787 , \comparator/n786 , \comparator/n785 ,
         \comparator/n784 , \comparator/n783 , \comparator/n782 ,
         \comparator/n781 , \comparator/n780 , \comparator/n779 ,
         \comparator/n778 , \comparator/n777 , \comparator/n776 ,
         \comparator/n775 , \comparator/n774 , \comparator/n773 ,
         \comparator/n772 , \comparator/n771 , \comparator/n770 ,
         \comparator/n769 , \comparator/n768 , \comparator/n767 ,
         \comparator/n766 , \comparator/n765 , \comparator/n764 ,
         \comparator/n763 , \comparator/n762 , \comparator/n761 ,
         \comparator/n760 , \comparator/n759 , \comparator/n758 ,
         \comparator/n757 , \comparator/n756 , \comparator/n755 ,
         \comparator/n754 , \comparator/n753 , \comparator/n752 ,
         \comparator/n751 , \comparator/n750 , \comparator/n749 ,
         \comparator/n748 , \comparator/n747 , \comparator/n746 ,
         \comparator/n745 , \comparator/n744 , \comparator/n743 ,
         \comparator/n742 , \comparator/n741 , \comparator/n740 ,
         \comparator/n739 , \comparator/n738 , \comparator/n737 ,
         \comparator/n736 , \comparator/n735 , \comparator/n734 ,
         \comparator/n733 , \comparator/n732 , \comparator/n731 ,
         \comparator/n730 , \comparator/n729 , \comparator/n728 ,
         \comparator/n727 , \comparator/n726 , \comparator/n725 ,
         \comparator/n724 , \comparator/n723 , \comparator/n722 ,
         \comparator/n721 , \comparator/n720 , \comparator/n719 ,
         \comparator/n718 , \comparator/n717 , \comparator/n716 ,
         \comparator/n715 , \comparator/n714 , \comparator/n713 ,
         \comparator/n712 , \comparator/n711 , \comparator/n710 ,
         \comparator/n709 , \comparator/n708 , \comparator/n707 ,
         \comparator/n706 , \comparator/n705 , \comparator/n704 ,
         \comparator/n703 , \comparator/n702 , \comparator/n701 ,
         \comparator/n700 , \comparator/n699 , \comparator/n698 ,
         \comparator/n697 , \comparator/n696 , \comparator/n695 ,
         \comparator/n694 , \comparator/n693 , \comparator/n692 ,
         \comparator/n691 , \comparator/n690 , \comparator/n689 ,
         \comparator/n688 , \comparator/n687 , \comparator/n686 ,
         \comparator/n685 , \comparator/n684 , \comparator/n683 ,
         \comparator/n682 , \comparator/n681 , \comparator/n680 ,
         \comparator/n679 , \comparator/n678 , \comparator/n677 ,
         \comparator/n676 , \comparator/n675 , \comparator/n674 ,
         \comparator/n673 , \comparator/n672 , \comparator/n671 ,
         \comparator/n670 , \comparator/n669 , \comparator/n668 ,
         \comparator/n667 , \comparator/n666 , \comparator/n665 ,
         \comparator/n664 , \comparator/n663 , \comparator/n662 ,
         \comparator/n661 , \comparator/n660 , \comparator/n659 ,
         \comparator/n658 , \comparator/n657 , \comparator/n656 ,
         \comparator/n655 , \comparator/n654 , \comparator/n653 ,
         \comparator/n652 , \comparator/n651 , \comparator/n650 ,
         \comparator/n649 , \comparator/n648 , \comparator/n647 ,
         \comparator/n646 , \comparator/n645 , \comparator/n644 ,
         \comparator/n643 , \comparator/n642 , \comparator/n641 ,
         \comparator/n640 , \comparator/n639 , \comparator/n638 ,
         \comparator/n637 , \comparator/n636 , \comparator/n635 ,
         \comparator/n634 , \comparator/n633 , \comparator/n632 ,
         \comparator/n631 , \comparator/n630 , \comparator/n629 ,
         \comparator/n628 , \comparator/n627 , \comparator/n626 ,
         \comparator/n625 , \comparator/n624 , \comparator/n623 ,
         \comparator/n622 , \comparator/n621 , \comparator/n620 ,
         \comparator/n619 , \comparator/n618 , \comparator/n617 ,
         \comparator/n616 , \comparator/n615 , \comparator/n614 ,
         \comparator/n613 , \comparator/n612 , \comparator/n611 ,
         \comparator/n610 , \comparator/n609 , \comparator/n608 ,
         \comparator/n607 , \comparator/n606 , \comparator/n605 ,
         \comparator/n604 , \comparator/n603 , \comparator/n602 ,
         \comparator/n601 , \comparator/n600 , \comparator/n599 ,
         \comparator/n598 , \comparator/n597 , \comparator/n596 ,
         \comparator/n595 , \comparator/n594 , \comparator/n593 ,
         \comparator/n592 , \comparator/n591 , \comparator/n590 ,
         \comparator/n589 , \comparator/n588 , \comparator/n587 ,
         \comparator/n586 , \comparator/n585 , \comparator/n584 ,
         \comparator/n583 , \comparator/n582 , \comparator/n581 ,
         \comparator/n580 , \comparator/n579 , \comparator/n578 ,
         \comparator/n577 , \comparator/n576 , \comparator/n575 ,
         \comparator/n574 , \comparator/n573 , \comparator/n572 ,
         \comparator/n571 , \comparator/n570 , \comparator/n569 ,
         \comparator/n568 , \comparator/n567 , \comparator/n566 ,
         \comparator/n565 , \comparator/n564 , \comparator/n563 ,
         \comparator/n562 , \comparator/n561 , \comparator/n560 ,
         \comparator/n559 , \comparator/n558 , \comparator/n557 ,
         \comparator/n556 , \comparator/n555 , \comparator/n554 ,
         \comparator/n553 , \comparator/n552 , \comparator/n551 ,
         \comparator/n550 , \comparator/n549 , \comparator/n548 ,
         \comparator/n547 , \comparator/n546 , \comparator/n545 ,
         \comparator/n544 , \comparator/n543 , \comparator/n542 ,
         \comparator/n541 , \comparator/n540 , \comparator/n539 ,
         \comparator/n538 , \comparator/n537 , \comparator/n536 ,
         \comparator/n535 , \comparator/n534 , \comparator/n533 ,
         \comparator/n532 , \comparator/n531 , \comparator/n530 ,
         \comparator/n529 , \comparator/n528 , \comparator/n527 ,
         \comparator/n526 , \comparator/n525 , \comparator/n524 ,
         \comparator/n523 , \comparator/n522 , \comparator/n521 ,
         \comparator/n520 , \comparator/n519 , \comparator/n518 ,
         \comparator/n517 , \comparator/n516 , \comparator/n515 ,
         \comparator/n514 , \comparator/n513 , \comparator/n512 ,
         \comparator/n511 , \comparator/n510 , \comparator/n509 ,
         \comparator/n508 , \comparator/n507 , \comparator/n506 ,
         \comparator/n505 , \comparator/n504 , \comparator/n503 ,
         \comparator/n502 , \comparator/n501 , \comparator/n500 ,
         \comparator/n499 , \comparator/n498 , \comparator/n497 ,
         \comparator/n496 , \comparator/n495 , \comparator/n494 ,
         \comparator/n493 , \comparator/n492 , \comparator/n491 ,
         \comparator/n490 , \comparator/n489 , \comparator/n488 ,
         \comparator/n487 , \comparator/n486 , \comparator/n485 ,
         \comparator/n484 , \comparator/n483 , \comparator/n482 ,
         \comparator/n481 , \comparator/n480 , \comparator/n479 ,
         \comparator/n478 , \comparator/n477 , \comparator/n476 ,
         \comparator/n475 , \comparator/n474 , \comparator/n473 ,
         \comparator/n472 , \comparator/n471 , \comparator/n470 ,
         \comparator/n469 , \comparator/n468 , \comparator/n467 ,
         \comparator/n466 , \comparator/n465 , \comparator/n464 ,
         \comparator/n463 , \comparator/n462 , \comparator/n461 ,
         \comparator/n460 , \comparator/n459 , \comparator/n458 ,
         \comparator/n457 , \comparator/n456 , \comparator/n455 ,
         \comparator/n454 , \comparator/n453 , \comparator/n452 ,
         \comparator/n451 , \comparator/n450 , \comparator/n449 ,
         \comparator/n448 , \comparator/n447 , \comparator/n446 ,
         \comparator/n445 , \comparator/n444 , \comparator/n443 ,
         \comparator/n442 , \comparator/n441 , \comparator/n440 ,
         \comparator/n439 , \comparator/n438 , \comparator/n437 ,
         \comparator/n436 , \comparator/n435 , \comparator/n434 ,
         \comparator/n433 , \comparator/n432 , \comparator/n431 ,
         \comparator/n430 , \comparator/n429 , \comparator/n428 ,
         \comparator/n427 , \comparator/n426 , \comparator/n425 ,
         \comparator/n424 , \comparator/n423 , \comparator/n422 ,
         \comparator/n421 , \comparator/n420 , \comparator/n419 ,
         \comparator/n418 , \comparator/n417 , \comparator/n416 ,
         \comparator/n415 , \comparator/n414 , \comparator/n413 ,
         \comparator/n412 , \comparator/n411 , \comparator/n410 ,
         \comparator/n409 , \comparator/n408 , \comparator/n407 ,
         \comparator/n406 , \comparator/n405 , \comparator/n404 ,
         \comparator/n403 , \comparator/n402 , \comparator/n401 ,
         \comparator/n400 , \comparator/n399 , \comparator/n398 ,
         \comparator/n397 , \comparator/n396 , \comparator/n395 ,
         \comparator/n394 , \comparator/n393 , \comparator/n392 ,
         \comparator/n391 , \comparator/n390 , \comparator/n389 ,
         \comparator/n388 , \comparator/n387 , \comparator/n386 ,
         \comparator/n385 , \comparator/n384 , \comparator/n383 ,
         \comparator/n382 , \comparator/n381 , \comparator/n380 ,
         \comparator/n379 , \comparator/n378 , \comparator/n377 ,
         \comparator/n376 , \comparator/n375 , \comparator/n374 ,
         \comparator/n373 , \comparator/n372 , \comparator/n371 ,
         \comparator/n370 , \comparator/n369 , \comparator/n368 ,
         \comparator/n367 , \comparator/n366 , \comparator/n365 ,
         \comparator/n364 , \comparator/n363 , \comparator/n362 ,
         \comparator/n361 , \comparator/n360 , \comparator/n359 ,
         \comparator/n358 , \comparator/n357 , \comparator/n356 ,
         \comparator/n355 , \comparator/n354 , \comparator/n353 ,
         \comparator/n352 , \comparator/n351 , \comparator/n350 ,
         \comparator/n349 , \comparator/n348 , \comparator/n347 ,
         \comparator/n346 , \comparator/n345 , \comparator/n344 ,
         \comparator/n343 , \comparator/n342 , \comparator/n341 ,
         \comparator/n340 , \comparator/n339 , \comparator/n338 ,
         \comparator/n337 , \comparator/n336 , \comparator/n335 ,
         \comparator/n334 , \comparator/n333 , \comparator/n332 ,
         \comparator/n331 , \comparator/n330 , \comparator/n329 ,
         \comparator/n328 , \comparator/n327 , \comparator/n326 ,
         \comparator/n325 , \comparator/n324 , \comparator/n323 ,
         \comparator/n322 , \comparator/n321 , \comparator/n320 ,
         \comparator/n319 , \comparator/n318 , \comparator/n317 ,
         \comparator/n316 , \comparator/n315 , \comparator/n314 ,
         \comparator/n313 , \comparator/n312 , \comparator/n311 ,
         \comparator/n310 , \comparator/n309 , \comparator/n308 ,
         \comparator/n307 , \comparator/n306 , \comparator/n305 ,
         \comparator/n304 , \comparator/n303 , \comparator/n302 ,
         \comparator/n301 , \comparator/n300 , \comparator/n299 ,
         \comparator/n298 , \comparator/n297 , \comparator/n296 ,
         \comparator/n295 , \comparator/n294 , \comparator/n293 ,
         \comparator/n292 , \comparator/n291 , \comparator/n290 ,
         \comparator/n289 , \comparator/n288 , \comparator/n287 ,
         \comparator/n286 , \comparator/n285 , \comparator/n284 ,
         \comparator/n283 , \comparator/n282 , \comparator/n281 ,
         \comparator/n280 , \comparator/n279 , \comparator/n278 ,
         \comparator/n277 , \comparator/n276 , \comparator/n275 ,
         \comparator/n274 , \comparator/n273 , \comparator/n272 ,
         \comparator/n271 , \comparator/n270 , \comparator/n269 ,
         \comparator/n268 , \comparator/n267 , \comparator/n266 ,
         \comparator/n265 , \comparator/n264 , \comparator/n263 ,
         \comparator/n262 , \comparator/n261 , \comparator/n260 ,
         \comparator/n259 , \comparator/n258 , \comparator/n257 ,
         \comparator/n256 , \comparator/n255 , \comparator/n254 ,
         \comparator/n253 , \comparator/n252 , \comparator/n251 ,
         \comparator/n250 , \comparator/n249 , \comparator/n248 ,
         \comparator/n247 , \comparator/n246 , \comparator/n245 ,
         \comparator/n244 , \comparator/n243 , \comparator/n242 ,
         \comparator/n241 , \comparator/n240 , \comparator/n239 ,
         \comparator/n238 , \comparator/n237 , \comparator/n236 ,
         \comparator/n235 , \comparator/n234 , \comparator/n233 ,
         \comparator/n232 , \comparator/n231 , \comparator/n230 ,
         \comparator/n229 , \comparator/n228 , \comparator/n227 ,
         \comparator/n226 , \comparator/n225 , \comparator/n224 ,
         \comparator/n223 , \comparator/n222 , \comparator/n221 ,
         \comparator/n220 , \comparator/n219 , \comparator/n218 ,
         \comparator/n217 , \comparator/n216 , \comparator/n215 ,
         \comparator/n214 , \comparator/n213 , \comparator/n212 ,
         \comparator/n211 , \comparator/n210 , \comparator/n209 ,
         \comparator/n208 , \comparator/n207 , \comparator/n206 ,
         \comparator/n205 , \comparator/n204 , \comparator/n203 ,
         \comparator/n202 , \comparator/n201 , \comparator/n200 ,
         \comparator/n199 , \comparator/n198 , \comparator/n197 ,
         \comparator/n196 , \comparator/n195 , \comparator/n194 ,
         \comparator/n193 , \comparator/n192 , \comparator/n191 ,
         \comparator/n190 , \comparator/n189 , \comparator/n188 ,
         \comparator/n187 , \comparator/n186 , \comparator/n185 ,
         \comparator/n184 , \comparator/n183 , \comparator/n182 ,
         \comparator/n181 , \comparator/n180 , \comparator/n179 ,
         \comparator/n178 , \comparator/n177 , \comparator/n176 ,
         \comparator/n175 , \comparator/n174 , \comparator/n173 ,
         \comparator/n172 , \comparator/n171 , \comparator/n170 ,
         \comparator/n169 , \comparator/n168 , \comparator/n167 ,
         \comparator/n166 , \comparator/n165 , \comparator/n164 ,
         \comparator/n163 , \comparator/n162 , \comparator/n161 ,
         \comparator/n160 , \comparator/n159 , \comparator/n158 ,
         \comparator/n157 , \comparator/n156 , \comparator/n155 ,
         \comparator/n154 , \comparator/n153 , \comparator/n152 ,
         \comparator/n151 , \comparator/n150 , \comparator/n149 ,
         \comparator/n148 , \comparator/n147 , \comparator/n146 ,
         \comparator/n145 , \comparator/n144 , \comparator/n143 ,
         \comparator/n142 , \comparator/n141 , \comparator/n140 ,
         \comparator/n139 , \comparator/n138 , \comparator/n137 ,
         \comparator/n136 , \comparator/n135 , \comparator/n134 ,
         \comparator/n133 , \comparator/n132 , \comparator/n131 ,
         \comparator/n130 , \comparator/n129 , \comparator/n128 ,
         \comparator/n127 , \comparator/n126 , \comparator/n125 ,
         \comparator/n124 , \comparator/n123 , \comparator/n122 ,
         \comparator/n121 , \comparator/n120 , \comparator/n119 ,
         \comparator/n118 , \comparator/n117 , \comparator/n116 ,
         \comparator/n115 , \comparator/n114 , \comparator/n113 ,
         \comparator/n112 , \comparator/n111 , \comparator/n110 ,
         \comparator/n109 , \comparator/n108 , \comparator/n107 ,
         \comparator/n106 , \comparator/n105 , \comparator/n104 ,
         \comparator/n103 , \comparator/n102 , \comparator/n101 ,
         \comparator/n100 , \comparator/n99 , \comparator/n98 ,
         \comparator/n97 , \comparator/n96 , \comparator/n95 ,
         \comparator/n94 , \comparator/n93 , \comparator/n92 ,
         \comparator/n91 , \comparator/n90 , \comparator/n89 ,
         \comparator/n88 , \comparator/n87 , \comparator/n86 ,
         \comparator/n85 , \comparator/n84 , \comparator/n83 ,
         \comparator/n82 , \comparator/n81 , \comparator/n80 ,
         \comparator/n79 , \comparator/n78 , \comparator/n77 ,
         \comparator/n76 , \comparator/n75 , \comparator/n74 ,
         \comparator/n73 , \comparator/n72 , \comparator/n71 ,
         \comparator/n70 , \comparator/n69 , \comparator/n68 ,
         \comparator/n67 , \comparator/n66 , \comparator/n65 ,
         \comparator/n64 , \comparator/n63 , \comparator/n62 ,
         \comparator/n61 , \comparator/n60 , \comparator/n59 ,
         \comparator/n58 , \comparator/n57 , \comparator/n56 ,
         \comparator/n55 , \comparator/n54 , \comparator/n53 ,
         \comparator/n52 , \comparator/n51 , \comparator/n50 ,
         \comparator/n49 , \comparator/n48 , \comparator/n47 ,
         \comparator/n46 , \comparator/n45 , \comparator/n44 ,
         \comparator/n43 , \comparator/n42 , \comparator/n41 ,
         \comparator/n40 , \comparator/n39 , \comparator/n38 ,
         \comparator/n37 , \comparator/n36 , \comparator/n35 ,
         \comparator/n34 , \comparator/n33 , \comparator/n32 ,
         \comparator/n31 , \comparator/n30 , \comparator/n29 ,
         \comparator/n28 , \comparator/n27 , \comparator/n26 ,
         \comparator/n25 , \comparator/n24 , \comparator/n23 ,
         \comparator/n22 , \comparator/n21 , \comparator/n20 ,
         \comparator/n19 , \comparator/n18 , \comparator/n17 ,
         \comparator/n16 , \comparator/n15 , \comparator/n14 ,
         \comparator/n13 , \comparator/n12 , \comparator/n11 ,
         \comparator/n10 , \comparator/n9 , \comparator/n8 , \comparator/n7 ,
         \comparator/n6 , \comparator/n5 , \comparator/n4 , \comparator/n3 ,
         \comparator/n2 , \comparator/n1 , \comparator/N2046 ,
         \comparator/N2045 , \comparator/N2044 , \comparator/N2043 ,
         \comparator/N2042 , \comparator/N2041 , \comparator/N2040 ,
         \comparator/N2039 , \comparator/N2038 , \comparator/N2037 ,
         \comparator/N2036 , \comparator/N2035 , \comparator/N2034 ,
         \comparator/N2033 , \comparator/N2032 , \comparator/N2031 ,
         \comparator/N2030 , \comparator/N2029 , \comparator/N2028 ,
         \comparator/N2027 , \comparator/N2026 , \comparator/N2025 ,
         \comparator/N2024 , \comparator/N2023 , \comparator/N2022 ,
         \comparator/N2021 , \comparator/N2020 , \comparator/N2019 ,
         \comparator/N2018 , \comparator/N2017 , \comparator/N2016 ,
         \comparator/N2015 , \comparator/N2014 , \comparator/N2013 ,
         \comparator/N2012 , \comparator/N2011 , \comparator/N2010 ,
         \comparator/N2009 , \comparator/N2008 , \comparator/N2007 ,
         \comparator/N2006 , \comparator/N2005 , \comparator/N2004 ,
         \comparator/N2003 , \comparator/N2002 , \comparator/N2001 ,
         \comparator/N2000 , \comparator/N1999 , \comparator/N1998 ,
         \comparator/N1997 , \comparator/N1996 , \comparator/N1995 ,
         \comparator/N1994 , \comparator/N1993 , \comparator/N1992 ,
         \comparator/N1991 , \comparator/N1990 , \comparator/N1989 ,
         \comparator/N1988 , \comparator/N1987 , \comparator/N1986 ,
         \comparator/N1985 , \comparator/N1984 , \comparator/N1983 ,
         \comparator/N1982 , \comparator/N1981 , \comparator/N1980 ,
         \comparator/N1979 , \comparator/N1978 , \comparator/N1977 ,
         \comparator/N1976 , \comparator/N1975 , \comparator/N1974 ,
         \comparator/N1973 , \comparator/N1972 , \comparator/N1971 ,
         \comparator/N1970 , \comparator/N1969 , \comparator/N1968 ,
         \comparator/N1967 , \comparator/N1966 , \comparator/N1965 ,
         \comparator/N1964 , \comparator/N1963 , \comparator/N1962 ,
         \comparator/N1961 , \comparator/N1960 , \comparator/N1959 ,
         \comparator/N1958 , \comparator/N1957 , \comparator/N1956 ,
         \comparator/N1955 , \comparator/N1954 , \comparator/N1953 ,
         \comparator/N1952 , \comparator/N1951 , \comparator/N1950 ,
         \comparator/N1949 , \comparator/N1948 , \comparator/N1947 ,
         \comparator/N1946 , \comparator/N1945 , \comparator/N1944 ,
         \comparator/N1943 , \comparator/N1942 , \comparator/N1941 ,
         \comparator/N1940 , \comparator/N1939 , \comparator/N1938 ,
         \comparator/N1937 , \comparator/N1936 , \comparator/N1935 ,
         \comparator/N1934 , \comparator/N1933 , \comparator/N1932 ,
         \comparator/N1931 , \comparator/N1930 , \comparator/N1929 ,
         \comparator/N1928 , \comparator/N1927 , \comparator/N1926 ,
         \comparator/N1925 , \comparator/N1924 , \comparator/N1923 ,
         \comparator/N1922 , \comparator/N1921 , \comparator/N1920 ,
         \comparator/N1919 , \comparator/N1918 , \comparator/N1917 ,
         \comparator/N1916 , \comparator/N1915 , \comparator/N1914 ,
         \comparator/N1913 , \comparator/N1912 , \comparator/N1911 ,
         \comparator/N1910 , \comparator/N1909 , \comparator/N1908 ,
         \comparator/N1907 , \comparator/N1906 , \comparator/N1905 ,
         \comparator/N1904 , \comparator/N1903 , \comparator/N1902 ,
         \comparator/N1901 , \comparator/N1900 , \comparator/N1899 ,
         \comparator/N1898 , \comparator/N1897 , \comparator/N1896 ,
         \comparator/N1895 , \comparator/N1894 , \comparator/N1893 ,
         \comparator/N1892 , \comparator/N1891 , \comparator/N1890 ,
         \comparator/N1889 , \comparator/N1888 , \comparator/N1887 ,
         \comparator/N1886 , \comparator/N1885 , \comparator/N1884 ,
         \comparator/N1883 , \comparator/N1882 , \comparator/N1881 ,
         \comparator/N1880 , \comparator/N1879 , \comparator/N1878 ,
         \comparator/N1877 , \comparator/N1876 , \comparator/N1875 ,
         \comparator/N1874 , \comparator/N1873 , \comparator/N1872 ,
         \comparator/N1871 , \comparator/N1870 , \comparator/N1869 ,
         \comparator/N1868 , \comparator/N1867 , \comparator/N1866 ,
         \comparator/N1865 , \comparator/N1864 , \comparator/N1863 ,
         \comparator/N1862 , \comparator/N1861 , \comparator/N1860 ,
         \comparator/N1859 , \comparator/N1858 , \comparator/N1857 ,
         \comparator/N1856 , \comparator/N1855 , \comparator/N1854 ,
         \comparator/N1853 , \comparator/N1852 , \comparator/N1851 ,
         \comparator/N1850 , \comparator/N1849 , \comparator/N1848 ,
         \comparator/N1847 , \comparator/N1846 , \comparator/N1845 ,
         \comparator/N1844 , \comparator/N1843 , \comparator/N1842 ,
         \comparator/N1841 , \comparator/N1840 , \comparator/N1839 ,
         \comparator/N1838 , \comparator/N1837 , \comparator/N1836 ,
         \comparator/N1835 , \comparator/N1834 , \comparator/N1833 ,
         \comparator/N1832 , \comparator/N1831 , \comparator/N1830 ,
         \comparator/N1829 , \comparator/N1828 , \comparator/N1827 ,
         \comparator/N1826 , \comparator/N1825 , \comparator/N1824 ,
         \comparator/N1823 , \comparator/N1822 , \comparator/N1821 ,
         \comparator/N1820 , \comparator/N1819 , \comparator/N1818 ,
         \comparator/N1817 , \comparator/N1816 , \comparator/N1815 ,
         \comparator/N1814 , \comparator/N1813 , \comparator/N1812 ,
         \comparator/N1811 , \comparator/N1810 , \comparator/N1809 ,
         \comparator/N1808 , \comparator/N1807 , \comparator/N1806 ,
         \comparator/N1805 , \comparator/N1804 , \comparator/N1803 ,
         \comparator/N1802 , \comparator/N1801 , \comparator/N1800 ,
         \comparator/N1799 , \comparator/N1798 , \comparator/N1797 ,
         \comparator/N1796 , \comparator/N1795 , \comparator/N1794 ,
         \comparator/N1793 , \comparator/N1792 , \comparator/N1791 ,
         \comparator/N1790 , \comparator/N1789 , \comparator/N1788 ,
         \comparator/N1787 , \comparator/N1786 , \comparator/N1785 ,
         \comparator/N1784 , \comparator/N1783 , \comparator/N1782 ,
         \comparator/N1781 , \comparator/N1780 , \comparator/N1779 ,
         \comparator/N1778 , \comparator/N1777 , \comparator/N1776 ,
         \comparator/N1775 , \comparator/N1774 , \comparator/N1773 ,
         \comparator/N1772 , \comparator/N1771 , \comparator/N1770 ,
         \comparator/N1769 , \comparator/N1768 , \comparator/N1767 ,
         \comparator/N1766 , \comparator/N1765 , \comparator/N1764 ,
         \comparator/N1763 , \comparator/N1762 , \comparator/N1761 ,
         \comparator/N1760 , \comparator/N1759 , \comparator/N1758 ,
         \comparator/N1757 , \comparator/N1756 , \comparator/N1755 ,
         \comparator/N1754 , \comparator/N1753 , \comparator/N1752 ,
         \comparator/N1751 , \comparator/N1750 , \comparator/N1749 ,
         \comparator/N1748 , \comparator/N1747 , \comparator/N1746 ,
         \comparator/N1745 , \comparator/N1744 , \comparator/N1743 ,
         \comparator/N1742 , \comparator/N1741 , \comparator/N1740 ,
         \comparator/N1739 , \comparator/N1738 , \comparator/N1737 ,
         \comparator/N1736 , \comparator/N1735 , \comparator/N1734 ,
         \comparator/N1733 , \comparator/N1732 , \comparator/N1731 ,
         \comparator/N1730 , \comparator/N1729 , \comparator/N1728 ,
         \comparator/N1727 , \comparator/N1726 , \comparator/N1725 ,
         \comparator/N1724 , \comparator/N1723 , \comparator/N1722 ,
         \comparator/N1721 , \comparator/N1720 , \comparator/N1719 ,
         \comparator/N1718 , \comparator/N1717 , \comparator/N1716 ,
         \comparator/N1715 , \comparator/N1714 , \comparator/N1713 ,
         \comparator/N1712 , \comparator/N1711 , \comparator/N1710 ,
         \comparator/N1709 , \comparator/N1708 , \comparator/N1707 ,
         \comparator/N1706 , \comparator/N1705 , \comparator/N1704 ,
         \comparator/N1703 , \comparator/N1702 , \comparator/N1701 ,
         \comparator/N1700 , \comparator/N1699 , \comparator/N1698 ,
         \comparator/N1697 , \comparator/N1696 , \comparator/N1695 ,
         \comparator/N1694 , \comparator/N1693 , \comparator/N1692 ,
         \comparator/N1691 , \comparator/N1690 , \comparator/N1689 ,
         \comparator/N1688 , \comparator/N1687 , \comparator/N1686 ,
         \comparator/N1685 , \comparator/N1684 , \comparator/N1683 ,
         \comparator/N1682 , \comparator/N1681 , \comparator/N1680 ,
         \comparator/N1679 , \comparator/N1678 , \comparator/N1677 ,
         \comparator/N1676 , \comparator/N1675 , \comparator/N1674 ,
         \comparator/N1673 , \comparator/N1672 , \comparator/N1671 ,
         \comparator/N1670 , \comparator/N1669 , \comparator/N1668 ,
         \comparator/N1667 , \comparator/N1666 , \comparator/N1665 ,
         \comparator/N1664 , \comparator/N1663 , \comparator/N1662 ,
         \comparator/N1661 , \comparator/N1660 , \comparator/N1659 ,
         \comparator/N1658 , \comparator/N1657 , \comparator/N1656 ,
         \comparator/N1655 , \comparator/N1654 , \comparator/N1653 ,
         \comparator/N1652 , \comparator/N1651 , \comparator/N1650 ,
         \comparator/N1649 , \comparator/N1648 , \comparator/N1647 ,
         \comparator/N1646 , \comparator/N1645 , \comparator/N1644 ,
         \comparator/N1643 , \comparator/N1642 , \comparator/N1641 ,
         \comparator/N1640 , \comparator/N1639 , \comparator/N1638 ,
         \comparator/N1637 , \comparator/N1636 , \comparator/N1635 ,
         \comparator/N1634 , \comparator/N1633 , \comparator/N1632 ,
         \comparator/N1631 , \comparator/N1630 , \comparator/N1629 ,
         \comparator/N1628 , \comparator/N1627 , \comparator/N1626 ,
         \comparator/N1625 , \comparator/N1624 , \comparator/N1623 ,
         \comparator/N1622 , \comparator/N1621 , \comparator/N1620 ,
         \comparator/N1619 , \comparator/N1618 , \comparator/N1617 ,
         \comparator/N1616 , \comparator/N1615 , \comparator/N1614 ,
         \comparator/N1613 , \comparator/N1612 , \comparator/N1611 ,
         \comparator/N1610 , \comparator/N1609 , \comparator/N1608 ,
         \comparator/N1607 , \comparator/N1606 , \comparator/N1605 ,
         \comparator/N1604 , \comparator/N1603 , \comparator/N1602 ,
         \comparator/N1601 , \comparator/N1600 , \comparator/N1599 ,
         \comparator/N1598 , \comparator/N1597 , \comparator/N1596 ,
         \comparator/N1595 , \comparator/N1594 , \comparator/N1593 ,
         \comparator/N1592 , \comparator/N1591 , \comparator/N1590 ,
         \comparator/N1589 , \comparator/N1588 , \comparator/N1587 ,
         \comparator/N1586 , \comparator/N1585 , \comparator/N1584 ,
         \comparator/N1583 , \comparator/N1582 , \comparator/N1581 ,
         \comparator/N1580 , \comparator/N1579 , \comparator/N1578 ,
         \comparator/N1577 , \comparator/N1576 , \comparator/N1575 ,
         \comparator/N1574 , \comparator/N1573 , \comparator/N1572 ,
         \comparator/N1571 , \comparator/N1570 , \comparator/N1569 ,
         \comparator/N1568 , \comparator/N1567 , \comparator/N1566 ,
         \comparator/N1565 , \comparator/N1564 , \comparator/N1563 ,
         \comparator/N1562 , \comparator/N1561 , \comparator/N1560 ,
         \comparator/N1559 , \comparator/N1558 , \comparator/N1557 ,
         \comparator/N1556 , \comparator/N1555 , \comparator/N1554 ,
         \comparator/N1553 , \comparator/N1552 , \comparator/N1551 ,
         \comparator/N1550 , \comparator/N1549 , \comparator/N1548 ,
         \comparator/N1547 , \comparator/N1546 , \comparator/N1545 ,
         \comparator/N1544 , \comparator/N1543 , \comparator/N1542 ,
         \comparator/N1541 , \comparator/N1540 , \comparator/N1539 ,
         \comparator/N1538 , \comparator/N1537 , \comparator/N1536 ,
         \comparator/N1535 , \comparator/N1534 , \comparator/N1533 ,
         \comparator/N1532 , \comparator/N1531 , \comparator/N1530 ,
         \comparator/N1529 , \comparator/N1528 , \comparator/N1527 ,
         \comparator/N1526 , \comparator/N1525 , \comparator/N1524 ,
         \comparator/N1523 , \comparator/N1522 , \comparator/N1521 ,
         \comparator/N1520 , \comparator/N1519 , \comparator/N1518 ,
         \comparator/N1517 , \comparator/N1516 , \comparator/N1515 ,
         \comparator/N1514 , \comparator/N1513 , \comparator/N1512 ,
         \comparator/N1511 , \comparator/N1510 , \comparator/N1509 ,
         \comparator/N1508 , \comparator/N1507 , \comparator/N1506 ,
         \comparator/N1505 , \comparator/N1504 , \comparator/N1503 ,
         \comparator/N1502 , \comparator/N1501 , \comparator/N1500 ,
         \comparator/N1499 , \comparator/N1498 , \comparator/N1497 ,
         \comparator/N1496 , \comparator/N1495 , \comparator/N1494 ,
         \comparator/N1493 , \comparator/N1492 , \comparator/N1491 ,
         \comparator/N1490 , \comparator/N1489 , \comparator/N1488 ,
         \comparator/N1487 , \comparator/N1486 , \comparator/N1485 ,
         \comparator/N1484 , \comparator/N1483 , \comparator/N1482 ,
         \comparator/N1481 , \comparator/N1480 , \comparator/N1479 ,
         \comparator/N1478 , \comparator/N1477 , \comparator/N1476 ,
         \comparator/N1475 , \comparator/N1474 , \comparator/N1473 ,
         \comparator/N1472 , \comparator/N1471 , \comparator/N1470 ,
         \comparator/N1469 , \comparator/N1468 , \comparator/N1467 ,
         \comparator/N1466 , \comparator/N1465 , \comparator/N1464 ,
         \comparator/N1463 , \comparator/N1462 , \comparator/N1461 ,
         \comparator/N1460 , \comparator/N1459 , \comparator/N1458 ,
         \comparator/N1457 , \comparator/N1456 , \comparator/N1455 ,
         \comparator/N1454 , \comparator/N1453 , \comparator/N1452 ,
         \comparator/N1451 , \comparator/N1450 , \comparator/N1449 ,
         \comparator/N1448 , \comparator/N1447 , \comparator/N1446 ,
         \comparator/N1445 , \comparator/N1444 , \comparator/N1443 ,
         \comparator/N1442 , \comparator/N1441 , \comparator/N1440 ,
         \comparator/N1439 , \comparator/N1438 , \comparator/N1437 ,
         \comparator/N1436 , \comparator/N1435 , \comparator/N1434 ,
         \comparator/N1433 , \comparator/N1432 , \comparator/N1431 ,
         \comparator/N1430 , \comparator/N1429 , \comparator/N1428 ,
         \comparator/N1427 , \comparator/N1426 , \comparator/N1425 ,
         \comparator/N1424 , \comparator/N1423 , \comparator/N1422 ,
         \comparator/N1421 , \comparator/N1420 , \comparator/N1419 ,
         \comparator/N1418 , \comparator/N1417 , \comparator/N1416 ,
         \comparator/N1415 , \comparator/N1414 , \comparator/N1413 ,
         \comparator/N1412 , \comparator/N1411 , \comparator/N1410 ,
         \comparator/N1409 , \comparator/N1408 , \comparator/N1407 ,
         \comparator/N1406 , \comparator/N1405 , \comparator/N1404 ,
         \comparator/N1403 , \comparator/N1402 , \comparator/N1401 ,
         \comparator/N1400 , \comparator/N1399 , \comparator/N1398 ,
         \comparator/N1397 , \comparator/N1396 , \comparator/N1395 ,
         \comparator/N1394 , \comparator/N1393 , \comparator/N1392 ,
         \comparator/N1391 , \comparator/N1390 , \comparator/N1389 ,
         \comparator/N1388 , \comparator/N1387 , \comparator/N1386 ,
         \comparator/N1385 , \comparator/N1384 , \comparator/N1383 ,
         \comparator/N1382 , \comparator/N1381 , \comparator/N1380 ,
         \comparator/N1379 , \comparator/N1378 , \comparator/N1377 ,
         \comparator/N1376 , \comparator/N1375 , \comparator/N1374 ,
         \comparator/N1373 , \comparator/N1372 , \comparator/N1371 ,
         \comparator/N1370 , \comparator/N1369 , \comparator/N1368 ,
         \comparator/N1367 , \comparator/N1366 , \comparator/N1365 ,
         \comparator/N1364 , \comparator/N1363 , \comparator/N1362 ,
         \comparator/N1361 , \comparator/N1360 , \comparator/N1359 ,
         \comparator/N1358 , \comparator/N1357 , \comparator/N1356 ,
         \comparator/N1355 , \comparator/N1354 , \comparator/N1353 ,
         \comparator/N1352 , \comparator/N1351 , \comparator/N1350 ,
         \comparator/N1349 , \comparator/N1348 , \comparator/N1347 ,
         \comparator/N1346 , \comparator/N1345 , \comparator/N1344 ,
         \comparator/N1343 , \comparator/N1342 , \comparator/N1341 ,
         \comparator/N1340 , \comparator/N1339 , \comparator/N1338 ,
         \comparator/N1337 , \comparator/N1336 , \comparator/N1335 ,
         \comparator/N1334 , \comparator/N1333 , \comparator/N1332 ,
         \comparator/N1331 , \comparator/N1330 , \comparator/N1329 ,
         \comparator/N1328 , \comparator/N1327 , \comparator/N1326 ,
         \comparator/N1325 , \comparator/N1324 , \comparator/N1323 ,
         \comparator/N1322 , \comparator/N1321 , \comparator/N1320 ,
         \comparator/N1319 , \comparator/N1318 , \comparator/N1317 ,
         \comparator/N1316 , \comparator/N1315 , \comparator/N1314 ,
         \comparator/N1313 , \comparator/N1312 , \comparator/N1311 ,
         \comparator/N1310 , \comparator/N1309 , \comparator/N1308 ,
         \comparator/N1307 , \comparator/N1306 , \comparator/N1305 ,
         \comparator/N1304 , \comparator/N1303 , \comparator/N1302 ,
         \comparator/N1301 , \comparator/N1300 , \comparator/N1299 ,
         \comparator/N1298 , \comparator/N1297 , \comparator/N1296 ,
         \comparator/N1295 , \comparator/N1294 , \comparator/N1293 ,
         \comparator/N1292 , \comparator/N1291 , \comparator/N1290 ,
         \comparator/N1289 , \comparator/N1288 , \comparator/N1287 ,
         \comparator/N1286 , \comparator/N1285 , \comparator/N1284 ,
         \comparator/N1283 , \comparator/N1282 , \comparator/N1281 ,
         \comparator/N1280 , \comparator/N1279 , \comparator/N1278 ,
         \comparator/N1277 , \comparator/N1276 , \comparator/N1275 ,
         \comparator/N1274 , \comparator/N1273 , \comparator/N1272 ,
         \comparator/N1271 , \comparator/N1270 , \comparator/N1269 ,
         \comparator/N1268 , \comparator/N1267 , \comparator/N1266 ,
         \comparator/N1265 , \comparator/N1264 , \comparator/N1263 ,
         \comparator/N1262 , \comparator/N1261 , \comparator/N1260 ,
         \comparator/N1259 , \comparator/N1258 , \comparator/N1257 ,
         \comparator/N1256 , \comparator/N1255 , \comparator/N1254 ,
         \comparator/N1253 , \comparator/N1252 , \comparator/N1251 ,
         \comparator/N1250 , \comparator/N1249 , \comparator/N1248 ,
         \comparator/N1247 , \comparator/N1246 , \comparator/N1245 ,
         \comparator/N1244 , \comparator/N1243 , \comparator/N1242 ,
         \comparator/N1241 , \comparator/N1240 , \comparator/N1239 ,
         \comparator/N1238 , \comparator/N1237 , \comparator/N1236 ,
         \comparator/N1235 , \comparator/N1234 , \comparator/N1233 ,
         \comparator/N1232 , \comparator/N1231 , \comparator/N1230 ,
         \comparator/N1229 , \comparator/N1228 , \comparator/N1227 ,
         \comparator/N1226 , \comparator/N1225 , \comparator/N1224 ,
         \comparator/N1223 , \comparator/N1222 , \comparator/N1221 ,
         \comparator/N1220 , \comparator/N1219 , \comparator/N1218 ,
         \comparator/N1217 , \comparator/N1216 , \comparator/N1215 ,
         \comparator/N1214 , \comparator/N1213 , \comparator/N1212 ,
         \comparator/N1211 , \comparator/N1210 , \comparator/N1209 ,
         \comparator/N1208 , \comparator/N1207 , \comparator/N1206 ,
         \comparator/N1205 , \comparator/N1204 , \comparator/N1203 ,
         \comparator/N1202 , \comparator/N1201 , \comparator/N1200 ,
         \comparator/N1199 , \comparator/N1198 , \comparator/N1197 ,
         \comparator/N1196 , \comparator/N1195 , \comparator/N1194 ,
         \comparator/N1193 , \comparator/N1192 , \comparator/N1191 ,
         \comparator/N1190 , \comparator/N1189 , \comparator/N1188 ,
         \comparator/N1187 , \comparator/N1186 , \comparator/N1185 ,
         \comparator/N1184 , \comparator/N1183 , \comparator/N1182 ,
         \comparator/N1181 , \comparator/N1180 , \comparator/N1179 ,
         \comparator/N1178 , \comparator/N1177 , \comparator/N1176 ,
         \comparator/N1175 , \comparator/N1174 , \comparator/N1173 ,
         \comparator/N1172 , \comparator/N1171 , \comparator/N1170 ,
         \comparator/N1169 , \comparator/N1168 , \comparator/N1167 ,
         \comparator/N1166 , \comparator/N1165 , \comparator/N1164 ,
         \comparator/N1163 , \comparator/N1162 , \comparator/N1161 ,
         \comparator/N1160 , \comparator/N1159 , \comparator/N1158 ,
         \comparator/N1157 , \comparator/N1156 , \comparator/N1155 ,
         \comparator/N1154 , \comparator/N1153 , \comparator/N1152 ,
         \comparator/N1151 , \comparator/N1150 , \comparator/N1149 ,
         \comparator/N1148 , \comparator/N1147 , \comparator/N1146 ,
         \comparator/N1145 , \comparator/N1144 , \comparator/N1143 ,
         \comparator/N1142 , \comparator/N1141 , \comparator/N1140 ,
         \comparator/N1139 , \comparator/N1138 , \comparator/N1137 ,
         \comparator/N1136 , \comparator/N1135 , \comparator/N1134 ,
         \comparator/N1133 , \comparator/N1132 , \comparator/N1131 ,
         \comparator/N1130 , \comparator/N1129 , \comparator/N1128 ,
         \comparator/N1127 , \comparator/N1126 , \comparator/N1125 ,
         \comparator/N1124 , \comparator/N1123 , \comparator/N1122 ,
         \comparator/N1121 , \comparator/N1120 , \comparator/N1119 ,
         \comparator/N1118 , \comparator/N1117 , \comparator/N1116 ,
         \comparator/N1115 , \comparator/N1114 , \comparator/N1113 ,
         \comparator/N1112 , \comparator/N1111 , \comparator/N1110 ,
         \comparator/N1109 , \comparator/N1108 , \comparator/N1107 ,
         \comparator/N1106 , \comparator/N1105 , \comparator/N1104 ,
         \comparator/N1103 , \comparator/N1102 , \comparator/N1101 ,
         \comparator/N1100 , \comparator/N1099 , \comparator/N1098 ,
         \comparator/N1097 , \comparator/N1096 , \comparator/N1095 ,
         \comparator/N1094 , \comparator/N1093 , \comparator/N1092 ,
         \comparator/N1091 , \comparator/N1090 , \comparator/N1089 ,
         \comparator/N1088 , \comparator/N1087 , \comparator/N1086 ,
         \comparator/N1085 , \comparator/N1084 , \comparator/N1083 ,
         \comparator/N1082 , \comparator/N1081 , \comparator/N1080 ,
         \comparator/N1079 , \comparator/N1078 , \comparator/N1077 ,
         \comparator/N1076 , \comparator/N1075 , \comparator/N1074 ,
         \comparator/N1073 , \comparator/N1072 , \comparator/N1071 ,
         \comparator/N1070 , \comparator/N1069 , \comparator/N1068 ,
         \comparator/N1067 , \comparator/N1066 , \comparator/N1065 ,
         \comparator/N1064 , \comparator/N1063 , \comparator/N1062 ,
         \comparator/N1061 , \comparator/N1060 , \comparator/N1059 ,
         \comparator/N1058 , \comparator/N1057 , \comparator/N1056 ,
         \comparator/N1055 , \comparator/N1054 , \comparator/N1053 ,
         \comparator/N1052 , \comparator/N1051 , \comparator/N1050 ,
         \comparator/N1049 , \comparator/N1048 , \comparator/N1047 ,
         \comparator/N1046 , \comparator/N1045 , \comparator/N1044 ,
         \comparator/N1043 , \comparator/N1042 , \comparator/N1041 ,
         \comparator/N1040 , \comparator/N1039 , \comparator/N1038 ,
         \comparator/N1037 , \comparator/N1036 , \comparator/N1035 ,
         \comparator/N1034 , \comparator/N1033 , \comparator/N1032 ,
         \comparator/N1031 , \comparator/N1030 , \comparator/N1029 ,
         \comparator/N1028 , \comparator/N1027 , \comparator/N1026 ,
         \comparator/N1025 , \comparator/N1024 , \comparator/N1023 ,
         \comparator/N1022 , \comparator/N1021 , \comparator/N1020 ,
         \comparator/N1019 , \comparator/N1018 , \comparator/N1017 ,
         \comparator/N1016 , \comparator/N1015 , \comparator/N1014 ,
         \comparator/N1013 , \comparator/N1012 , \comparator/N1011 ,
         \comparator/N1010 , \comparator/N1009 , \comparator/N1008 ,
         \comparator/N1007 , \comparator/N1006 , \comparator/N1005 ,
         \comparator/N1004 , \comparator/N1003 , \comparator/N1002 ,
         \comparator/N1001 , \comparator/N1000 , \comparator/N999 ,
         \comparator/N998 , \comparator/N997 , \comparator/N996 ,
         \comparator/N995 , \comparator/N994 , \comparator/N993 ,
         \comparator/N992 , \comparator/N991 , \comparator/N990 ,
         \comparator/N989 , \comparator/N988 , \comparator/N987 ,
         \comparator/N986 , \comparator/N985 , \comparator/N984 ,
         \comparator/N983 , \comparator/N982 , \comparator/N981 ,
         \comparator/N980 , \comparator/N979 , \comparator/N978 ,
         \comparator/N977 , \comparator/N976 , \comparator/N975 ,
         \comparator/N974 , \comparator/N973 , \comparator/N972 ,
         \comparator/N971 , \comparator/N970 , \comparator/N969 ,
         \comparator/N968 , \comparator/N967 , \comparator/N966 ,
         \comparator/N965 , \comparator/N964 , \comparator/N963 ,
         \comparator/N962 , \comparator/N961 , \comparator/N960 ,
         \comparator/N959 , \comparator/N958 , \comparator/N957 ,
         \comparator/N956 , \comparator/N955 , \comparator/N954 ,
         \comparator/N953 , \comparator/N952 , \comparator/N951 ,
         \comparator/N950 , \comparator/N949 , \comparator/N948 ,
         \comparator/N947 , \comparator/N946 , \comparator/N945 ,
         \comparator/N944 , \comparator/N943 , \comparator/N942 ,
         \comparator/N941 , \comparator/N940 , \comparator/N939 ,
         \comparator/N938 , \comparator/N937 , \comparator/N936 ,
         \comparator/N935 , \comparator/N934 , \comparator/N933 ,
         \comparator/N932 , \comparator/N931 , \comparator/N930 ,
         \comparator/N929 , \comparator/N928 , \comparator/N927 ,
         \comparator/N926 , \comparator/N925 , \comparator/N924 ,
         \comparator/N923 , \comparator/N922 , \comparator/N921 ,
         \comparator/N920 , \comparator/N919 , \comparator/N918 ,
         \comparator/N917 , \comparator/N916 , \comparator/N915 ,
         \comparator/N914 , \comparator/N913 , \comparator/N912 ,
         \comparator/N911 , \comparator/N910 , \comparator/N909 ,
         \comparator/N908 , \comparator/N907 , \comparator/N906 ,
         \comparator/N905 , \comparator/N904 , \comparator/N903 ,
         \comparator/N902 , \comparator/N901 , \comparator/N900 ,
         \comparator/N899 , \comparator/N898 , \comparator/N897 ,
         \comparator/N896 , \comparator/N895 , \comparator/N894 ,
         \comparator/N893 , \comparator/N892 , \comparator/N891 ,
         \comparator/N890 , \comparator/N889 , \comparator/N888 ,
         \comparator/N887 , \comparator/N886 , \comparator/N885 ,
         \comparator/N884 , \comparator/N883 , \comparator/N882 ,
         \comparator/N881 , \comparator/N880 , \comparator/N879 ,
         \comparator/N878 , \comparator/N877 , \comparator/N876 ,
         \comparator/N875 , \comparator/N874 , \comparator/N873 ,
         \comparator/N872 , \comparator/N871 , \comparator/N870 ,
         \comparator/N869 , \comparator/N868 , \comparator/N867 ,
         \comparator/N866 , \comparator/N865 , \comparator/N864 ,
         \comparator/N863 , \comparator/N862 , \comparator/N861 ,
         \comparator/N860 , \comparator/N859 , \comparator/N858 ,
         \comparator/N857 , \comparator/N856 , \comparator/N855 ,
         \comparator/N854 , \comparator/N853 , \comparator/N852 ,
         \comparator/N851 , \comparator/N850 , \comparator/N849 ,
         \comparator/N848 , \comparator/N847 , \comparator/N846 ,
         \comparator/N845 , \comparator/N844 , \comparator/N843 ,
         \comparator/N842 , \comparator/N841 , \comparator/N840 ,
         \comparator/N839 , \comparator/N838 , \comparator/N837 ,
         \comparator/N836 , \comparator/N835 , \comparator/N834 ,
         \comparator/N833 , \comparator/N832 , \comparator/N831 ,
         \comparator/N830 , \comparator/N829 , \comparator/N828 ,
         \comparator/N827 , \comparator/N826 , \comparator/N825 ,
         \comparator/N824 , \comparator/N823 , \comparator/N822 ,
         \comparator/N821 , \comparator/N820 , \comparator/N819 ,
         \comparator/N818 , \comparator/N817 , \comparator/N816 ,
         \comparator/N815 , \comparator/N814 , \comparator/N813 ,
         \comparator/N812 , \comparator/N811 , \comparator/N810 ,
         \comparator/N809 , \comparator/N808 , \comparator/N807 ,
         \comparator/N806 , \comparator/N805 , \comparator/N804 ,
         \comparator/N803 , \comparator/N802 , \comparator/N801 ,
         \comparator/N800 , \comparator/N799 , \comparator/N798 ,
         \comparator/N797 , \comparator/N796 , \comparator/N795 ,
         \comparator/N794 , \comparator/N793 , \comparator/N792 ,
         \comparator/N791 , \comparator/N790 , \comparator/N789 ,
         \comparator/N788 , \comparator/N787 , \comparator/N786 ,
         \comparator/N785 , \comparator/N784 , \comparator/N783 ,
         \comparator/N782 , \comparator/N781 , \comparator/N780 ,
         \comparator/N779 , \comparator/N778 , \comparator/N777 ,
         \comparator/N776 , \comparator/N775 , \comparator/N774 ,
         \comparator/N773 , \comparator/N772 , \comparator/N771 ,
         \comparator/N770 , \comparator/N769 , \comparator/N768 ,
         \comparator/N767 , \comparator/N766 , \comparator/N765 ,
         \comparator/N764 , \comparator/N763 , \comparator/N762 ,
         \comparator/N761 , \comparator/N760 , \comparator/N759 ,
         \comparator/N758 , \comparator/N757 , \comparator/N756 ,
         \comparator/N755 , \comparator/N754 , \comparator/N753 ,
         \comparator/N752 , \comparator/N751 , \comparator/N750 ,
         \comparator/N749 , \comparator/N748 , \comparator/N747 ,
         \comparator/N746 , \comparator/N745 , \comparator/N744 ,
         \comparator/N743 , \comparator/N742 , \comparator/N741 ,
         \comparator/N740 , \comparator/N739 , \comparator/N738 ,
         \comparator/N737 , \comparator/N736 , \comparator/N735 ,
         \comparator/N734 , \comparator/N733 , \comparator/N732 ,
         \comparator/N731 , \comparator/N730 , \comparator/N729 ,
         \comparator/N728 , \comparator/N727 , \comparator/N726 ,
         \comparator/N725 , \comparator/N724 , \comparator/N723 ,
         \comparator/N722 , \comparator/N721 , \comparator/N720 ,
         \comparator/N719 , \comparator/N718 , \comparator/N717 ,
         \comparator/N716 , \comparator/N715 , \comparator/N714 ,
         \comparator/N713 , \comparator/N712 , \comparator/N711 ,
         \comparator/N710 , \comparator/N709 , \comparator/N708 ,
         \comparator/N707 , \comparator/N706 , \comparator/N705 ,
         \comparator/N704 , \comparator/N703 , \comparator/N702 ,
         \comparator/N701 , \comparator/N700 , \comparator/N699 ,
         \comparator/N698 , \comparator/N697 , \comparator/N696 ,
         \comparator/N695 , \comparator/N694 , \comparator/N693 ,
         \comparator/N692 , \comparator/N691 , \comparator/N690 ,
         \comparator/N689 , \comparator/N688 , \comparator/N687 ,
         \comparator/N686 , \comparator/N685 , \comparator/N684 ,
         \comparator/N683 , \comparator/N682 , \comparator/N681 ,
         \comparator/N680 , \comparator/N679 , \comparator/N678 ,
         \comparator/N677 , \comparator/N676 , \comparator/N675 ,
         \comparator/N674 , \comparator/N673 , \comparator/N672 ,
         \comparator/N671 , \comparator/N670 , \comparator/N669 ,
         \comparator/N668 , \comparator/N667 , \comparator/N666 ,
         \comparator/N665 , \comparator/N664 , \comparator/N663 ,
         \comparator/N662 , \comparator/N661 , \comparator/N660 ,
         \comparator/N659 , \comparator/N658 , \comparator/N657 ,
         \comparator/N656 , \comparator/N655 , \comparator/N654 ,
         \comparator/N653 , \comparator/N652 , \comparator/N651 ,
         \comparator/N650 , \comparator/N649 , \comparator/N648 ,
         \comparator/N647 , \comparator/N646 , \comparator/N645 ,
         \comparator/N644 , \comparator/N643 , \comparator/N642 ,
         \comparator/N641 , \comparator/N640 , \comparator/N639 ,
         \comparator/N638 , \comparator/N637 , \comparator/N636 ,
         \comparator/N635 , \comparator/N634 , \comparator/N633 ,
         \comparator/N632 , \comparator/N631 , \comparator/N630 ,
         \comparator/N629 , \comparator/N628 , \comparator/N627 ,
         \comparator/N626 , \comparator/N625 , \comparator/N624 ,
         \comparator/N623 , \comparator/N622 , \comparator/N621 ,
         \comparator/N620 , \comparator/N619 , \comparator/N618 ,
         \comparator/N617 , \comparator/N616 , \comparator/N615 ,
         \comparator/N614 , \comparator/N613 , \comparator/N612 ,
         \comparator/N611 , \comparator/N610 , \comparator/N609 ,
         \comparator/N608 , \comparator/N607 , \comparator/N606 ,
         \comparator/N605 , \comparator/N604 , \comparator/N603 ,
         \comparator/N602 , \comparator/N601 , \comparator/N600 ,
         \comparator/N599 , \comparator/N598 , \comparator/N597 ,
         \comparator/N596 , \comparator/N595 , \comparator/N594 ,
         \comparator/N593 , \comparator/N592 , \comparator/N591 ,
         \comparator/N590 , \comparator/N589 , \comparator/N588 ,
         \comparator/N587 , \comparator/N586 , \comparator/N585 ,
         \comparator/N584 , \comparator/N583 , \comparator/N582 ,
         \comparator/N581 , \comparator/N580 , \comparator/N579 ,
         \comparator/N578 , \comparator/N577 , \comparator/N576 ,
         \comparator/N575 , \comparator/N574 , \comparator/N573 ,
         \comparator/N572 , \comparator/N571 , \comparator/N570 ,
         \comparator/N569 , \comparator/N568 , \comparator/N567 ,
         \comparator/N566 , \comparator/N565 , \comparator/N564 ,
         \comparator/N563 , \comparator/N562 , \comparator/N561 ,
         \comparator/N560 , \comparator/N559 , \comparator/N558 ,
         \comparator/N557 , \comparator/N556 , \comparator/N555 ,
         \comparator/N554 , \comparator/N553 , \comparator/N552 ,
         \comparator/N551 , \comparator/N550 , \comparator/N549 ,
         \comparator/N548 , \comparator/N547 , \comparator/N546 ,
         \comparator/N545 , \comparator/N544 , \comparator/N543 ,
         \comparator/N542 , \comparator/N541 , \comparator/N540 ,
         \comparator/N539 , \comparator/N538 , \comparator/N537 ,
         \comparator/N536 , \comparator/N535 , \comparator/N534 ,
         \comparator/N533 , \comparator/N532 , \comparator/N531 ,
         \comparator/N530 , \comparator/N529 , \comparator/N528 ,
         \comparator/N527 , \comparator/N526 , \comparator/N525 ,
         \comparator/N524 , \comparator/N523 , \comparator/N522 ,
         \comparator/N521 , \comparator/N520 , \comparator/N519 ,
         \comparator/N518 , \comparator/N517 , \comparator/N516 ,
         \comparator/N515 , \comparator/N514 , \comparator/N513 ,
         \comparator/N512 , \comparator/N511 , \comparator/N510 ,
         \comparator/N509 , \comparator/N508 , \comparator/N507 ,
         \comparator/N506 , \comparator/N505 , \comparator/N504 ,
         \comparator/N503 , \comparator/N502 , \comparator/N501 ,
         \comparator/N500 , \comparator/N499 , \comparator/N498 ,
         \comparator/N497 , \comparator/N496 , \comparator/N495 ,
         \comparator/N494 , \comparator/N493 , \comparator/N492 ,
         \comparator/N491 , \comparator/N490 , \comparator/N489 ,
         \comparator/N488 , \comparator/N487 , \comparator/N486 ,
         \comparator/N485 , \comparator/N484 , \comparator/N483 ,
         \comparator/N482 , \comparator/N481 , \comparator/N480 ,
         \comparator/N479 , \comparator/N478 , \comparator/N477 ,
         \comparator/N476 , \comparator/N475 , \comparator/N474 ,
         \comparator/N473 , \comparator/N472 , \comparator/N471 ,
         \comparator/N470 , \comparator/N469 , \comparator/N468 ,
         \comparator/N467 , \comparator/N466 , \comparator/N465 ,
         \comparator/N464 , \comparator/N463 , \comparator/N462 ,
         \comparator/N461 , \comparator/N460 , \comparator/N459 ,
         \comparator/N458 , \comparator/N457 , \comparator/N456 ,
         \comparator/N455 , \comparator/N454 , \comparator/N453 ,
         \comparator/N452 , \comparator/N451 , \comparator/N450 ,
         \comparator/N449 , \comparator/N448 , \comparator/N447 ,
         \comparator/N446 , \comparator/N445 , \comparator/N444 ,
         \comparator/N443 , \comparator/N442 , \comparator/N441 ,
         \comparator/N440 , \comparator/N439 , \comparator/N438 ,
         \comparator/N437 , \comparator/N436 , \comparator/N435 ,
         \comparator/N434 , \comparator/N433 , \comparator/N432 ,
         \comparator/N431 , \comparator/N430 , \comparator/N429 ,
         \comparator/N428 , \comparator/N427 , \comparator/N426 ,
         \comparator/N425 , \comparator/N424 , \comparator/N423 ,
         \comparator/N422 , \comparator/N421 , \comparator/N420 ,
         \comparator/N419 , \comparator/N418 , \comparator/N417 ,
         \comparator/N416 , \comparator/N415 , \comparator/N414 ,
         \comparator/N413 , \comparator/N412 , \comparator/N411 ,
         \comparator/N410 , \comparator/N409 , \comparator/N408 ,
         \comparator/N407 , \comparator/N406 , \comparator/N405 ,
         \comparator/N404 , \comparator/N403 , \comparator/N402 ,
         \comparator/N401 , \comparator/N400 , \comparator/N399 ,
         \comparator/N398 , \comparator/N397 , \comparator/N396 ,
         \comparator/N395 , \comparator/N394 , \comparator/N393 ,
         \comparator/N392 , \comparator/N391 , \comparator/N390 ,
         \comparator/N389 , \comparator/N388 , \comparator/N387 ,
         \comparator/N386 , \comparator/N385 , \comparator/N384 ,
         \comparator/N383 , \comparator/N382 , \comparator/N381 ,
         \comparator/N380 , \comparator/N379 , \comparator/N378 ,
         \comparator/N377 , \comparator/N376 , \comparator/N375 ,
         \comparator/N374 , \comparator/N373 , \comparator/N372 ,
         \comparator/N371 , \comparator/N370 , \comparator/N369 ,
         \comparator/N368 , \comparator/N367 , \comparator/N366 ,
         \comparator/N365 , \comparator/N364 , \comparator/N363 ,
         \comparator/N362 , \comparator/N361 , \comparator/N360 ,
         \comparator/N359 , \comparator/N358 , \comparator/N357 ,
         \comparator/N356 , \comparator/N355 , \comparator/N354 ,
         \comparator/N353 , \comparator/N352 , \comparator/N351 ,
         \comparator/N350 , \comparator/N349 , \comparator/N348 ,
         \comparator/N347 , \comparator/N346 , \comparator/N345 ,
         \comparator/N344 , \comparator/N343 , \comparator/N342 ,
         \comparator/N341 , \comparator/N340 , \comparator/N339 ,
         \comparator/N338 , \comparator/N337 , \comparator/N336 ,
         \comparator/N335 , \comparator/N334 , \comparator/N333 ,
         \comparator/N332 , \comparator/N331 , \comparator/N330 ,
         \comparator/N329 , \comparator/N328 , \comparator/N327 ,
         \comparator/N326 , \comparator/N325 , \comparator/N324 ,
         \comparator/N323 , \comparator/N322 , \comparator/N321 ,
         \comparator/N320 , \comparator/N319 , \comparator/N318 ,
         \comparator/N317 , \comparator/N316 , \comparator/N315 ,
         \comparator/N314 , \comparator/N313 , \comparator/N312 ,
         \comparator/N311 , \comparator/N310 , \comparator/N309 ,
         \comparator/N308 , \comparator/N307 , \comparator/N306 ,
         \comparator/N305 , \comparator/N304 , \comparator/N303 ,
         \comparator/N302 , \comparator/N301 , \comparator/N300 ,
         \comparator/N299 , \comparator/N298 , \comparator/N297 ,
         \comparator/N296 , \comparator/N295 , \comparator/N294 ,
         \comparator/N293 , \comparator/N292 , \comparator/N291 ,
         \comparator/N290 , \comparator/N289 , \comparator/N288 ,
         \comparator/N287 , \comparator/N286 , \comparator/N285 ,
         \comparator/N284 , \comparator/N283 , \comparator/N282 ,
         \comparator/N281 , \comparator/N280 , \comparator/N279 ,
         \comparator/N278 , \comparator/N277 , \comparator/N276 ,
         \comparator/N275 , \comparator/N274 , \comparator/N273 ,
         \comparator/N272 , \comparator/N271 , \comparator/N270 ,
         \comparator/N269 , \comparator/N268 , \comparator/N267 ,
         \comparator/N266 , \comparator/N265 , \comparator/N264 ,
         \comparator/N263 , \comparator/N262 , \comparator/N261 ,
         \comparator/N260 , \comparator/N259 , \comparator/N258 ,
         \comparator/N257 , \comparator/N256 , \comparator/N255 ,
         \comparator/N254 , \comparator/N253 , \comparator/N252 ,
         \comparator/N251 , \comparator/N250 , \comparator/N249 ,
         \comparator/N248 , \comparator/N247 , \comparator/N246 ,
         \comparator/N245 , \comparator/N244 , \comparator/N243 ,
         \comparator/N242 , \comparator/N241 , \comparator/N240 ,
         \comparator/N239 , \comparator/N238 , \comparator/N237 ,
         \comparator/N236 , \comparator/N235 , \comparator/N234 ,
         \comparator/N233 , \comparator/N232 , \comparator/N231 ,
         \comparator/N230 , \comparator/N229 , \comparator/N228 ,
         \comparator/N227 , \comparator/N226 , \comparator/N225 ,
         \comparator/N224 , \comparator/N223 , \comparator/N222 ,
         \comparator/N221 , \comparator/N220 , \comparator/N219 ,
         \comparator/N218 , \comparator/N217 , \comparator/N216 ,
         \comparator/N215 , \comparator/N214 , \comparator/N213 ,
         \comparator/N212 , \comparator/N211 , \comparator/N210 ,
         \comparator/N209 , \comparator/N208 , \comparator/N207 ,
         \comparator/N206 , \comparator/N205 , \comparator/N204 ,
         \comparator/N203 , \comparator/N202 , \comparator/N201 ,
         \comparator/N200 , \comparator/N199 , \comparator/N198 ,
         \comparator/N197 , \comparator/N196 , \comparator/N195 ,
         \comparator/N194 , \comparator/N193 , \comparator/N192 ,
         \comparator/N191 , \comparator/N190 , \comparator/N189 ,
         \comparator/N188 , \comparator/N187 , \comparator/N186 ,
         \comparator/N185 , \comparator/N184 , \comparator/N183 ,
         \comparator/N182 , \comparator/N181 , \comparator/N180 ,
         \comparator/N179 , \comparator/N178 , \comparator/N177 ,
         \comparator/N176 , \comparator/N175 , \comparator/N174 ,
         \comparator/N173 , \comparator/N172 , \comparator/N171 ,
         \comparator/N170 , \comparator/N169 , \comparator/N168 ,
         \comparator/N167 , \comparator/N166 , \comparator/N165 ,
         \comparator/N164 , \comparator/N163 , \comparator/N162 ,
         \comparator/N161 , \comparator/N160 , \comparator/N159 ,
         \comparator/N158 , \comparator/N157 , \comparator/N156 ,
         \comparator/N155 , \comparator/N154 , \comparator/N153 ,
         \comparator/N152 , \comparator/N151 , \comparator/N150 ,
         \comparator/N149 , \comparator/N148 , \comparator/N147 ,
         \comparator/N146 , \comparator/N145 , \comparator/N144 ,
         \comparator/N143 , \comparator/N142 , \comparator/N141 ,
         \comparator/N140 , \comparator/N139 , \comparator/N138 ,
         \comparator/N137 , \comparator/N136 , \comparator/N135 ,
         \comparator/N134 , \comparator/N133 , \comparator/N132 ,
         \comparator/N131 , \comparator/N130 , \comparator/N129 ,
         \comparator/N128 , \comparator/N127 , \comparator/N126 ,
         \comparator/N125 , \comparator/N124 , \comparator/N123 ,
         \comparator/N122 , \comparator/N121 , \comparator/N120 ,
         \comparator/N119 , \comparator/N118 , \comparator/N117 ,
         \comparator/N116 , \comparator/N115 , \comparator/N114 ,
         \comparator/N113 , \comparator/N112 , \comparator/N111 ,
         \comparator/N110 , \comparator/N109 , \comparator/N108 ,
         \comparator/N107 , \comparator/N106 , \comparator/N105 ,
         \comparator/N104 , \comparator/N103 , \comparator/N102 ,
         \comparator/N101 , \comparator/N100 , \comparator/N99 ,
         \comparator/N98 , \comparator/N97 , \comparator/N96 ,
         \comparator/N95 , \comparator/N94 , \comparator/N93 ,
         \comparator/N92 , \comparator/N91 , \comparator/N90 ,
         \comparator/N89 , \comparator/N88 , \comparator/N87 ,
         \comparator/N86 , \comparator/N85 , \comparator/N84 ,
         \comparator/N83 , \comparator/N82 , \comparator/N81 ,
         \comparator/N80 , \comparator/N79 , \comparator/N78 ,
         \comparator/N77 , \comparator/N76 , \comparator/N75 ,
         \comparator/N74 , \comparator/N73 , \comparator/N72 ,
         \comparator/N71 , \comparator/N70 , \comparator/N69 ,
         \comparator/N68 , \comparator/N67 , \comparator/N66 ,
         \comparator/N65 , \comparator/N64 , \comparator/N63 ,
         \comparator/N62 , \comparator/N61 , \comparator/N60 ,
         \comparator/N59 , \comparator/N58 , \comparator/N57 ,
         \comparator/N56 , \comparator/N55 , \comparator/N54 ,
         \comparator/N53 , \comparator/N52 , \comparator/N51 ,
         \comparator/N50 , \comparator/N49 , \comparator/N48 ,
         \comparator/N47 , \comparator/N46 , \comparator/N45 ,
         \comparator/N44 , \comparator/N43 , \comparator/N42 ,
         \comparator/N41 , \comparator/N40 , \comparator/N39 ,
         \comparator/N38 , \comparator/N37 , \comparator/N36 ,
         \comparator/N35 , \comparator/N34 , \comparator/N33 ,
         \comparator/N32 , \comparator/N31 , \comparator/N30 ,
         \comparator/N29 , \comparator/N28 , \comparator/N27 ,
         \comparator/N26 , \comparator/N25 , \comparator/N24 ,
         \comparator/N23 , \comparator/N22 , \comparator/N21 ,
         \comparator/N20 , \comparator/N19 , \comparator/N18 ,
         \comparator/N17 , \comparator/N16 , \comparator/N15 ,
         \comparator/N14 , \comparator/N13 , \comparator/N12 ,
         \comparator/N11 , \comparator/N10 , \comparator/N9 , \comparator/N8 ,
         \comparator/N7 , \comparator/N6 , \comparator/N5 , \comparator/N4 ,
         \comparator/N3 , \comparator/N2 , \comparator/N1 , \comparator/N0 ,
         \sig_prgm_register/clear_not , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  wire   [1023:0] a;
  wire   [1023:0] b;
  wire   [1023:0] \prgm_register/or_signal ;
  wire   [1023:0] \sig_prgm_register/or_signal ;

  inv \prgm_register/I_0  ( .a(clr), .out(\prgm_register/clear_not ) );
  inv \prgm_register/I_1  ( .a(enable), .out(\prgm_register/en_not ) );
  nand2 \prgm_register/C3082  ( .a(enable), .b(prgm), .out(\prgm_register/n1 )
         );
  nand2 \prgm_register/C3083  ( .a(\prgm_register/en_not ), .b(a[0]), .out(
        \prgm_register/n2 ) );
  nand2 \prgm_register/C3084  ( .a(\prgm_register/n1 ), .b(\prgm_register/n2 ), 
        .out(\prgm_register/or_signal [0]) );
  nand2 \prgm_register/C3085  ( .a(enable), .b(a[0]), .out(\prgm_register/n3 )
         );
  nand2 \prgm_register/C3086  ( .a(\prgm_register/en_not ), .b(a[1]), .out(
        \prgm_register/n4 ) );
  nand2 \prgm_register/C3087  ( .a(\prgm_register/n3 ), .b(\prgm_register/n4 ), 
        .out(\prgm_register/or_signal [1]) );
  nand2 \prgm_register/C3088  ( .a(enable), .b(a[1]), .out(\prgm_register/n5 )
         );
  nand2 \prgm_register/C3089  ( .a(\prgm_register/en_not ), .b(a[2]), .out(
        \prgm_register/n6 ) );
  nand2 \prgm_register/C3090  ( .a(\prgm_register/n5 ), .b(\prgm_register/n6 ), 
        .out(\prgm_register/or_signal [2]) );
  nand2 \prgm_register/C3091  ( .a(enable), .b(a[2]), .out(\prgm_register/n7 )
         );
  nand2 \prgm_register/C3092  ( .a(\prgm_register/en_not ), .b(a[3]), .out(
        \prgm_register/n8 ) );
  nand2 \prgm_register/C3093  ( .a(\prgm_register/n7 ), .b(\prgm_register/n8 ), 
        .out(\prgm_register/or_signal [3]) );
  nand2 \prgm_register/C3094  ( .a(enable), .b(a[3]), .out(\prgm_register/n9 )
         );
  nand2 \prgm_register/C3095  ( .a(\prgm_register/en_not ), .b(a[4]), .out(
        \prgm_register/n10 ) );
  nand2 \prgm_register/C3096  ( .a(\prgm_register/n9 ), .b(\prgm_register/n10 ), .out(\prgm_register/or_signal [4]) );
  nand2 \prgm_register/C3097  ( .a(enable), .b(a[4]), .out(\prgm_register/n11 ) );
  nand2 \prgm_register/C3098  ( .a(\prgm_register/en_not ), .b(a[5]), .out(
        \prgm_register/n12 ) );
  nand2 \prgm_register/C3099  ( .a(\prgm_register/n11 ), .b(
        \prgm_register/n12 ), .out(\prgm_register/or_signal [5]) );
  nand2 \prgm_register/C3100  ( .a(enable), .b(a[5]), .out(\prgm_register/n13 ) );
  nand2 \prgm_register/C3101  ( .a(\prgm_register/en_not ), .b(a[6]), .out(
        \prgm_register/n14 ) );
  nand2 \prgm_register/C3102  ( .a(\prgm_register/n13 ), .b(
        \prgm_register/n14 ), .out(\prgm_register/or_signal [6]) );
  nand2 \prgm_register/C3103  ( .a(enable), .b(a[6]), .out(\prgm_register/n15 ) );
  nand2 \prgm_register/C3104  ( .a(\prgm_register/en_not ), .b(a[7]), .out(
        \prgm_register/n16 ) );
  nand2 \prgm_register/C3105  ( .a(\prgm_register/n15 ), .b(
        \prgm_register/n16 ), .out(\prgm_register/or_signal [7]) );
  nand2 \prgm_register/C3106  ( .a(enable), .b(a[7]), .out(\prgm_register/n17 ) );
  nand2 \prgm_register/C3107  ( .a(\prgm_register/en_not ), .b(a[8]), .out(
        \prgm_register/n18 ) );
  nand2 \prgm_register/C3108  ( .a(\prgm_register/n17 ), .b(
        \prgm_register/n18 ), .out(\prgm_register/or_signal [8]) );
  nand2 \prgm_register/C3109  ( .a(enable), .b(a[8]), .out(\prgm_register/n19 ) );
  nand2 \prgm_register/C3110  ( .a(\prgm_register/en_not ), .b(a[9]), .out(
        \prgm_register/n20 ) );
  nand2 \prgm_register/C3111  ( .a(\prgm_register/n19 ), .b(
        \prgm_register/n20 ), .out(\prgm_register/or_signal [9]) );
  nand2 \prgm_register/C3112  ( .a(enable), .b(a[9]), .out(\prgm_register/n21 ) );
  nand2 \prgm_register/C3113  ( .a(\prgm_register/en_not ), .b(a[10]), .out(
        \prgm_register/n22 ) );
  nand2 \prgm_register/C3114  ( .a(\prgm_register/n21 ), .b(
        \prgm_register/n22 ), .out(\prgm_register/or_signal [10]) );
  nand2 \prgm_register/C3115  ( .a(enable), .b(a[10]), .out(
        \prgm_register/n23 ) );
  nand2 \prgm_register/C3116  ( .a(\prgm_register/en_not ), .b(a[11]), .out(
        \prgm_register/n24 ) );
  nand2 \prgm_register/C3117  ( .a(\prgm_register/n23 ), .b(
        \prgm_register/n24 ), .out(\prgm_register/or_signal [11]) );
  nand2 \prgm_register/C3118  ( .a(enable), .b(a[11]), .out(
        \prgm_register/n25 ) );
  nand2 \prgm_register/C3119  ( .a(\prgm_register/en_not ), .b(a[12]), .out(
        \prgm_register/n26 ) );
  nand2 \prgm_register/C3120  ( .a(\prgm_register/n25 ), .b(
        \prgm_register/n26 ), .out(\prgm_register/or_signal [12]) );
  nand2 \prgm_register/C3121  ( .a(enable), .b(a[12]), .out(
        \prgm_register/n27 ) );
  nand2 \prgm_register/C3122  ( .a(\prgm_register/en_not ), .b(a[13]), .out(
        \prgm_register/n28 ) );
  nand2 \prgm_register/C3123  ( .a(\prgm_register/n27 ), .b(
        \prgm_register/n28 ), .out(\prgm_register/or_signal [13]) );
  nand2 \prgm_register/C3124  ( .a(enable), .b(a[13]), .out(
        \prgm_register/n29 ) );
  nand2 \prgm_register/C3125  ( .a(\prgm_register/en_not ), .b(a[14]), .out(
        \prgm_register/n30 ) );
  nand2 \prgm_register/C3126  ( .a(\prgm_register/n29 ), .b(
        \prgm_register/n30 ), .out(\prgm_register/or_signal [14]) );
  nand2 \prgm_register/C3127  ( .a(enable), .b(a[14]), .out(
        \prgm_register/n31 ) );
  nand2 \prgm_register/C3128  ( .a(\prgm_register/en_not ), .b(a[15]), .out(
        \prgm_register/n32 ) );
  nand2 \prgm_register/C3129  ( .a(\prgm_register/n31 ), .b(
        \prgm_register/n32 ), .out(\prgm_register/or_signal [15]) );
  nand2 \prgm_register/C3130  ( .a(enable), .b(a[15]), .out(
        \prgm_register/n33 ) );
  nand2 \prgm_register/C3131  ( .a(\prgm_register/en_not ), .b(a[16]), .out(
        \prgm_register/n34 ) );
  nand2 \prgm_register/C3132  ( .a(\prgm_register/n33 ), .b(
        \prgm_register/n34 ), .out(\prgm_register/or_signal [16]) );
  nand2 \prgm_register/C3133  ( .a(enable), .b(a[16]), .out(
        \prgm_register/n35 ) );
  nand2 \prgm_register/C3134  ( .a(\prgm_register/en_not ), .b(a[17]), .out(
        \prgm_register/n36 ) );
  nand2 \prgm_register/C3135  ( .a(\prgm_register/n35 ), .b(
        \prgm_register/n36 ), .out(\prgm_register/or_signal [17]) );
  nand2 \prgm_register/C3136  ( .a(enable), .b(a[17]), .out(
        \prgm_register/n37 ) );
  nand2 \prgm_register/C3137  ( .a(\prgm_register/en_not ), .b(a[18]), .out(
        \prgm_register/n38 ) );
  nand2 \prgm_register/C3138  ( .a(\prgm_register/n37 ), .b(
        \prgm_register/n38 ), .out(\prgm_register/or_signal [18]) );
  nand2 \prgm_register/C3139  ( .a(enable), .b(a[18]), .out(
        \prgm_register/n39 ) );
  nand2 \prgm_register/C3140  ( .a(\prgm_register/en_not ), .b(a[19]), .out(
        \prgm_register/n40 ) );
  nand2 \prgm_register/C3141  ( .a(\prgm_register/n39 ), .b(
        \prgm_register/n40 ), .out(\prgm_register/or_signal [19]) );
  nand2 \prgm_register/C3142  ( .a(enable), .b(a[19]), .out(
        \prgm_register/n41 ) );
  nand2 \prgm_register/C3143  ( .a(\prgm_register/en_not ), .b(a[20]), .out(
        \prgm_register/n42 ) );
  nand2 \prgm_register/C3144  ( .a(\prgm_register/n41 ), .b(
        \prgm_register/n42 ), .out(\prgm_register/or_signal [20]) );
  nand2 \prgm_register/C3145  ( .a(enable), .b(a[20]), .out(
        \prgm_register/n43 ) );
  nand2 \prgm_register/C3146  ( .a(\prgm_register/en_not ), .b(a[21]), .out(
        \prgm_register/n44 ) );
  nand2 \prgm_register/C3147  ( .a(\prgm_register/n43 ), .b(
        \prgm_register/n44 ), .out(\prgm_register/or_signal [21]) );
  nand2 \prgm_register/C3148  ( .a(enable), .b(a[21]), .out(
        \prgm_register/n45 ) );
  nand2 \prgm_register/C3149  ( .a(\prgm_register/en_not ), .b(a[22]), .out(
        \prgm_register/n46 ) );
  nand2 \prgm_register/C3150  ( .a(\prgm_register/n45 ), .b(
        \prgm_register/n46 ), .out(\prgm_register/or_signal [22]) );
  nand2 \prgm_register/C3151  ( .a(enable), .b(a[22]), .out(
        \prgm_register/n47 ) );
  nand2 \prgm_register/C3152  ( .a(\prgm_register/en_not ), .b(a[23]), .out(
        \prgm_register/n48 ) );
  nand2 \prgm_register/C3153  ( .a(\prgm_register/n47 ), .b(
        \prgm_register/n48 ), .out(\prgm_register/or_signal [23]) );
  nand2 \prgm_register/C3154  ( .a(enable), .b(a[23]), .out(
        \prgm_register/n49 ) );
  nand2 \prgm_register/C3155  ( .a(\prgm_register/en_not ), .b(a[24]), .out(
        \prgm_register/n50 ) );
  nand2 \prgm_register/C3156  ( .a(\prgm_register/n49 ), .b(
        \prgm_register/n50 ), .out(\prgm_register/or_signal [24]) );
  nand2 \prgm_register/C3157  ( .a(enable), .b(a[24]), .out(
        \prgm_register/n51 ) );
  nand2 \prgm_register/C3158  ( .a(\prgm_register/en_not ), .b(a[25]), .out(
        \prgm_register/n52 ) );
  nand2 \prgm_register/C3159  ( .a(\prgm_register/n51 ), .b(
        \prgm_register/n52 ), .out(\prgm_register/or_signal [25]) );
  nand2 \prgm_register/C3160  ( .a(enable), .b(a[25]), .out(
        \prgm_register/n53 ) );
  nand2 \prgm_register/C3161  ( .a(\prgm_register/en_not ), .b(a[26]), .out(
        \prgm_register/n54 ) );
  nand2 \prgm_register/C3162  ( .a(\prgm_register/n53 ), .b(
        \prgm_register/n54 ), .out(\prgm_register/or_signal [26]) );
  nand2 \prgm_register/C3163  ( .a(enable), .b(a[26]), .out(
        \prgm_register/n55 ) );
  nand2 \prgm_register/C3164  ( .a(\prgm_register/en_not ), .b(a[27]), .out(
        \prgm_register/n56 ) );
  nand2 \prgm_register/C3165  ( .a(\prgm_register/n55 ), .b(
        \prgm_register/n56 ), .out(\prgm_register/or_signal [27]) );
  nand2 \prgm_register/C3166  ( .a(enable), .b(a[27]), .out(
        \prgm_register/n57 ) );
  nand2 \prgm_register/C3167  ( .a(\prgm_register/en_not ), .b(a[28]), .out(
        \prgm_register/n58 ) );
  nand2 \prgm_register/C3168  ( .a(\prgm_register/n57 ), .b(
        \prgm_register/n58 ), .out(\prgm_register/or_signal [28]) );
  nand2 \prgm_register/C3169  ( .a(enable), .b(a[28]), .out(
        \prgm_register/n59 ) );
  nand2 \prgm_register/C3170  ( .a(\prgm_register/en_not ), .b(a[29]), .out(
        \prgm_register/n60 ) );
  nand2 \prgm_register/C3171  ( .a(\prgm_register/n59 ), .b(
        \prgm_register/n60 ), .out(\prgm_register/or_signal [29]) );
  nand2 \prgm_register/C3172  ( .a(enable), .b(a[29]), .out(
        \prgm_register/n61 ) );
  nand2 \prgm_register/C3173  ( .a(\prgm_register/en_not ), .b(a[30]), .out(
        \prgm_register/n62 ) );
  nand2 \prgm_register/C3174  ( .a(\prgm_register/n61 ), .b(
        \prgm_register/n62 ), .out(\prgm_register/or_signal [30]) );
  nand2 \prgm_register/C3175  ( .a(enable), .b(a[30]), .out(
        \prgm_register/n63 ) );
  nand2 \prgm_register/C3176  ( .a(\prgm_register/en_not ), .b(a[31]), .out(
        \prgm_register/n64 ) );
  nand2 \prgm_register/C3177  ( .a(\prgm_register/n63 ), .b(
        \prgm_register/n64 ), .out(\prgm_register/or_signal [31]) );
  nand2 \prgm_register/C3178  ( .a(enable), .b(a[31]), .out(
        \prgm_register/n65 ) );
  nand2 \prgm_register/C3179  ( .a(\prgm_register/en_not ), .b(a[32]), .out(
        \prgm_register/n66 ) );
  nand2 \prgm_register/C3180  ( .a(\prgm_register/n65 ), .b(
        \prgm_register/n66 ), .out(\prgm_register/or_signal [32]) );
  nand2 \prgm_register/C3181  ( .a(enable), .b(a[32]), .out(
        \prgm_register/n67 ) );
  nand2 \prgm_register/C3182  ( .a(\prgm_register/en_not ), .b(a[33]), .out(
        \prgm_register/n68 ) );
  nand2 \prgm_register/C3183  ( .a(\prgm_register/n67 ), .b(
        \prgm_register/n68 ), .out(\prgm_register/or_signal [33]) );
  nand2 \prgm_register/C3184  ( .a(enable), .b(a[33]), .out(
        \prgm_register/n69 ) );
  nand2 \prgm_register/C3185  ( .a(\prgm_register/en_not ), .b(a[34]), .out(
        \prgm_register/n70 ) );
  nand2 \prgm_register/C3186  ( .a(\prgm_register/n69 ), .b(
        \prgm_register/n70 ), .out(\prgm_register/or_signal [34]) );
  nand2 \prgm_register/C3187  ( .a(enable), .b(a[34]), .out(
        \prgm_register/n71 ) );
  nand2 \prgm_register/C3188  ( .a(\prgm_register/en_not ), .b(a[35]), .out(
        \prgm_register/n72 ) );
  nand2 \prgm_register/C3189  ( .a(\prgm_register/n71 ), .b(
        \prgm_register/n72 ), .out(\prgm_register/or_signal [35]) );
  nand2 \prgm_register/C3190  ( .a(enable), .b(a[35]), .out(
        \prgm_register/n73 ) );
  nand2 \prgm_register/C3191  ( .a(\prgm_register/en_not ), .b(a[36]), .out(
        \prgm_register/n74 ) );
  nand2 \prgm_register/C3192  ( .a(\prgm_register/n73 ), .b(
        \prgm_register/n74 ), .out(\prgm_register/or_signal [36]) );
  nand2 \prgm_register/C3193  ( .a(enable), .b(a[36]), .out(
        \prgm_register/n75 ) );
  nand2 \prgm_register/C3194  ( .a(\prgm_register/en_not ), .b(a[37]), .out(
        \prgm_register/n76 ) );
  nand2 \prgm_register/C3195  ( .a(\prgm_register/n75 ), .b(
        \prgm_register/n76 ), .out(\prgm_register/or_signal [37]) );
  nand2 \prgm_register/C3196  ( .a(enable), .b(a[37]), .out(
        \prgm_register/n77 ) );
  nand2 \prgm_register/C3197  ( .a(\prgm_register/en_not ), .b(a[38]), .out(
        \prgm_register/n78 ) );
  nand2 \prgm_register/C3198  ( .a(\prgm_register/n77 ), .b(
        \prgm_register/n78 ), .out(\prgm_register/or_signal [38]) );
  nand2 \prgm_register/C3199  ( .a(enable), .b(a[38]), .out(
        \prgm_register/n79 ) );
  nand2 \prgm_register/C3200  ( .a(\prgm_register/en_not ), .b(a[39]), .out(
        \prgm_register/n80 ) );
  nand2 \prgm_register/C3201  ( .a(\prgm_register/n79 ), .b(
        \prgm_register/n80 ), .out(\prgm_register/or_signal [39]) );
  nand2 \prgm_register/C3202  ( .a(enable), .b(a[39]), .out(
        \prgm_register/n81 ) );
  nand2 \prgm_register/C3203  ( .a(\prgm_register/en_not ), .b(a[40]), .out(
        \prgm_register/n82 ) );
  nand2 \prgm_register/C3204  ( .a(\prgm_register/n81 ), .b(
        \prgm_register/n82 ), .out(\prgm_register/or_signal [40]) );
  nand2 \prgm_register/C3205  ( .a(enable), .b(a[40]), .out(
        \prgm_register/n83 ) );
  nand2 \prgm_register/C3206  ( .a(\prgm_register/en_not ), .b(a[41]), .out(
        \prgm_register/n84 ) );
  nand2 \prgm_register/C3207  ( .a(\prgm_register/n83 ), .b(
        \prgm_register/n84 ), .out(\prgm_register/or_signal [41]) );
  nand2 \prgm_register/C3208  ( .a(enable), .b(a[41]), .out(
        \prgm_register/n85 ) );
  nand2 \prgm_register/C3209  ( .a(\prgm_register/en_not ), .b(a[42]), .out(
        \prgm_register/n86 ) );
  nand2 \prgm_register/C3210  ( .a(\prgm_register/n85 ), .b(
        \prgm_register/n86 ), .out(\prgm_register/or_signal [42]) );
  nand2 \prgm_register/C3211  ( .a(enable), .b(a[42]), .out(
        \prgm_register/n87 ) );
  nand2 \prgm_register/C3212  ( .a(\prgm_register/en_not ), .b(a[43]), .out(
        \prgm_register/n88 ) );
  nand2 \prgm_register/C3213  ( .a(\prgm_register/n87 ), .b(
        \prgm_register/n88 ), .out(\prgm_register/or_signal [43]) );
  nand2 \prgm_register/C3214  ( .a(enable), .b(a[43]), .out(
        \prgm_register/n89 ) );
  nand2 \prgm_register/C3215  ( .a(\prgm_register/en_not ), .b(a[44]), .out(
        \prgm_register/n90 ) );
  nand2 \prgm_register/C3216  ( .a(\prgm_register/n89 ), .b(
        \prgm_register/n90 ), .out(\prgm_register/or_signal [44]) );
  nand2 \prgm_register/C3217  ( .a(enable), .b(a[44]), .out(
        \prgm_register/n91 ) );
  nand2 \prgm_register/C3218  ( .a(\prgm_register/en_not ), .b(a[45]), .out(
        \prgm_register/n92 ) );
  nand2 \prgm_register/C3219  ( .a(\prgm_register/n91 ), .b(
        \prgm_register/n92 ), .out(\prgm_register/or_signal [45]) );
  nand2 \prgm_register/C3220  ( .a(enable), .b(a[45]), .out(
        \prgm_register/n93 ) );
  nand2 \prgm_register/C3221  ( .a(\prgm_register/en_not ), .b(a[46]), .out(
        \prgm_register/n94 ) );
  nand2 \prgm_register/C3222  ( .a(\prgm_register/n93 ), .b(
        \prgm_register/n94 ), .out(\prgm_register/or_signal [46]) );
  nand2 \prgm_register/C3223  ( .a(enable), .b(a[46]), .out(
        \prgm_register/n95 ) );
  nand2 \prgm_register/C3224  ( .a(\prgm_register/en_not ), .b(a[47]), .out(
        \prgm_register/n96 ) );
  nand2 \prgm_register/C3225  ( .a(\prgm_register/n95 ), .b(
        \prgm_register/n96 ), .out(\prgm_register/or_signal [47]) );
  nand2 \prgm_register/C3226  ( .a(enable), .b(a[47]), .out(
        \prgm_register/n97 ) );
  nand2 \prgm_register/C3227  ( .a(\prgm_register/en_not ), .b(a[48]), .out(
        \prgm_register/n98 ) );
  nand2 \prgm_register/C3228  ( .a(\prgm_register/n97 ), .b(
        \prgm_register/n98 ), .out(\prgm_register/or_signal [48]) );
  nand2 \prgm_register/C3229  ( .a(enable), .b(a[48]), .out(
        \prgm_register/n99 ) );
  nand2 \prgm_register/C3230  ( .a(\prgm_register/en_not ), .b(a[49]), .out(
        \prgm_register/n100 ) );
  nand2 \prgm_register/C3231  ( .a(\prgm_register/n99 ), .b(
        \prgm_register/n100 ), .out(\prgm_register/or_signal [49]) );
  nand2 \prgm_register/C3232  ( .a(enable), .b(a[49]), .out(
        \prgm_register/n101 ) );
  nand2 \prgm_register/C3233  ( .a(\prgm_register/en_not ), .b(a[50]), .out(
        \prgm_register/n102 ) );
  nand2 \prgm_register/C3234  ( .a(\prgm_register/n101 ), .b(
        \prgm_register/n102 ), .out(\prgm_register/or_signal [50]) );
  nand2 \prgm_register/C3235  ( .a(enable), .b(a[50]), .out(
        \prgm_register/n103 ) );
  nand2 \prgm_register/C3236  ( .a(\prgm_register/en_not ), .b(a[51]), .out(
        \prgm_register/n104 ) );
  nand2 \prgm_register/C3237  ( .a(\prgm_register/n103 ), .b(
        \prgm_register/n104 ), .out(\prgm_register/or_signal [51]) );
  nand2 \prgm_register/C3238  ( .a(enable), .b(a[51]), .out(
        \prgm_register/n105 ) );
  nand2 \prgm_register/C3239  ( .a(\prgm_register/en_not ), .b(a[52]), .out(
        \prgm_register/n106 ) );
  nand2 \prgm_register/C3240  ( .a(\prgm_register/n105 ), .b(
        \prgm_register/n106 ), .out(\prgm_register/or_signal [52]) );
  nand2 \prgm_register/C3241  ( .a(enable), .b(a[52]), .out(
        \prgm_register/n107 ) );
  nand2 \prgm_register/C3242  ( .a(\prgm_register/en_not ), .b(a[53]), .out(
        \prgm_register/n108 ) );
  nand2 \prgm_register/C3243  ( .a(\prgm_register/n107 ), .b(
        \prgm_register/n108 ), .out(\prgm_register/or_signal [53]) );
  nand2 \prgm_register/C3244  ( .a(enable), .b(a[53]), .out(
        \prgm_register/n109 ) );
  nand2 \prgm_register/C3245  ( .a(\prgm_register/en_not ), .b(a[54]), .out(
        \prgm_register/n110 ) );
  nand2 \prgm_register/C3246  ( .a(\prgm_register/n109 ), .b(
        \prgm_register/n110 ), .out(\prgm_register/or_signal [54]) );
  nand2 \prgm_register/C3247  ( .a(enable), .b(a[54]), .out(
        \prgm_register/n111 ) );
  nand2 \prgm_register/C3248  ( .a(\prgm_register/en_not ), .b(a[55]), .out(
        \prgm_register/n112 ) );
  nand2 \prgm_register/C3249  ( .a(\prgm_register/n111 ), .b(
        \prgm_register/n112 ), .out(\prgm_register/or_signal [55]) );
  nand2 \prgm_register/C3250  ( .a(enable), .b(a[55]), .out(
        \prgm_register/n113 ) );
  nand2 \prgm_register/C3251  ( .a(\prgm_register/en_not ), .b(a[56]), .out(
        \prgm_register/n114 ) );
  nand2 \prgm_register/C3252  ( .a(\prgm_register/n113 ), .b(
        \prgm_register/n114 ), .out(\prgm_register/or_signal [56]) );
  nand2 \prgm_register/C3253  ( .a(enable), .b(a[56]), .out(
        \prgm_register/n115 ) );
  nand2 \prgm_register/C3254  ( .a(\prgm_register/en_not ), .b(a[57]), .out(
        \prgm_register/n116 ) );
  nand2 \prgm_register/C3255  ( .a(\prgm_register/n115 ), .b(
        \prgm_register/n116 ), .out(\prgm_register/or_signal [57]) );
  nand2 \prgm_register/C3256  ( .a(enable), .b(a[57]), .out(
        \prgm_register/n117 ) );
  nand2 \prgm_register/C3257  ( .a(\prgm_register/en_not ), .b(a[58]), .out(
        \prgm_register/n118 ) );
  nand2 \prgm_register/C3258  ( .a(\prgm_register/n117 ), .b(
        \prgm_register/n118 ), .out(\prgm_register/or_signal [58]) );
  nand2 \prgm_register/C3259  ( .a(enable), .b(a[58]), .out(
        \prgm_register/n119 ) );
  nand2 \prgm_register/C3260  ( .a(\prgm_register/en_not ), .b(a[59]), .out(
        \prgm_register/n120 ) );
  nand2 \prgm_register/C3261  ( .a(\prgm_register/n119 ), .b(
        \prgm_register/n120 ), .out(\prgm_register/or_signal [59]) );
  nand2 \prgm_register/C3262  ( .a(enable), .b(a[59]), .out(
        \prgm_register/n121 ) );
  nand2 \prgm_register/C3263  ( .a(\prgm_register/en_not ), .b(a[60]), .out(
        \prgm_register/n122 ) );
  nand2 \prgm_register/C3264  ( .a(\prgm_register/n121 ), .b(
        \prgm_register/n122 ), .out(\prgm_register/or_signal [60]) );
  nand2 \prgm_register/C3265  ( .a(enable), .b(a[60]), .out(
        \prgm_register/n123 ) );
  nand2 \prgm_register/C3266  ( .a(\prgm_register/en_not ), .b(a[61]), .out(
        \prgm_register/n124 ) );
  nand2 \prgm_register/C3267  ( .a(\prgm_register/n123 ), .b(
        \prgm_register/n124 ), .out(\prgm_register/or_signal [61]) );
  nand2 \prgm_register/C3268  ( .a(enable), .b(a[61]), .out(
        \prgm_register/n125 ) );
  nand2 \prgm_register/C3269  ( .a(\prgm_register/en_not ), .b(a[62]), .out(
        \prgm_register/n126 ) );
  nand2 \prgm_register/C3270  ( .a(\prgm_register/n125 ), .b(
        \prgm_register/n126 ), .out(\prgm_register/or_signal [62]) );
  nand2 \prgm_register/C3271  ( .a(enable), .b(a[62]), .out(
        \prgm_register/n127 ) );
  nand2 \prgm_register/C3272  ( .a(\prgm_register/en_not ), .b(a[63]), .out(
        \prgm_register/n128 ) );
  nand2 \prgm_register/C3273  ( .a(\prgm_register/n127 ), .b(
        \prgm_register/n128 ), .out(\prgm_register/or_signal [63]) );
  nand2 \prgm_register/C3274  ( .a(enable), .b(a[63]), .out(
        \prgm_register/n129 ) );
  nand2 \prgm_register/C3275  ( .a(\prgm_register/en_not ), .b(a[64]), .out(
        \prgm_register/n130 ) );
  nand2 \prgm_register/C3276  ( .a(\prgm_register/n129 ), .b(
        \prgm_register/n130 ), .out(\prgm_register/or_signal [64]) );
  nand2 \prgm_register/C3277  ( .a(enable), .b(a[64]), .out(
        \prgm_register/n131 ) );
  nand2 \prgm_register/C3278  ( .a(\prgm_register/en_not ), .b(a[65]), .out(
        \prgm_register/n132 ) );
  nand2 \prgm_register/C3279  ( .a(\prgm_register/n131 ), .b(
        \prgm_register/n132 ), .out(\prgm_register/or_signal [65]) );
  nand2 \prgm_register/C3280  ( .a(enable), .b(a[65]), .out(
        \prgm_register/n133 ) );
  nand2 \prgm_register/C3281  ( .a(\prgm_register/en_not ), .b(a[66]), .out(
        \prgm_register/n134 ) );
  nand2 \prgm_register/C3282  ( .a(\prgm_register/n133 ), .b(
        \prgm_register/n134 ), .out(\prgm_register/or_signal [66]) );
  nand2 \prgm_register/C3283  ( .a(enable), .b(a[66]), .out(
        \prgm_register/n135 ) );
  nand2 \prgm_register/C3284  ( .a(\prgm_register/en_not ), .b(a[67]), .out(
        \prgm_register/n136 ) );
  nand2 \prgm_register/C3285  ( .a(\prgm_register/n135 ), .b(
        \prgm_register/n136 ), .out(\prgm_register/or_signal [67]) );
  nand2 \prgm_register/C3286  ( .a(enable), .b(a[67]), .out(
        \prgm_register/n137 ) );
  nand2 \prgm_register/C3287  ( .a(\prgm_register/en_not ), .b(a[68]), .out(
        \prgm_register/n138 ) );
  nand2 \prgm_register/C3288  ( .a(\prgm_register/n137 ), .b(
        \prgm_register/n138 ), .out(\prgm_register/or_signal [68]) );
  nand2 \prgm_register/C3289  ( .a(enable), .b(a[68]), .out(
        \prgm_register/n139 ) );
  nand2 \prgm_register/C3290  ( .a(\prgm_register/en_not ), .b(a[69]), .out(
        \prgm_register/n140 ) );
  nand2 \prgm_register/C3291  ( .a(\prgm_register/n139 ), .b(
        \prgm_register/n140 ), .out(\prgm_register/or_signal [69]) );
  nand2 \prgm_register/C3292  ( .a(enable), .b(a[69]), .out(
        \prgm_register/n141 ) );
  nand2 \prgm_register/C3293  ( .a(\prgm_register/en_not ), .b(a[70]), .out(
        \prgm_register/n142 ) );
  nand2 \prgm_register/C3294  ( .a(\prgm_register/n141 ), .b(
        \prgm_register/n142 ), .out(\prgm_register/or_signal [70]) );
  nand2 \prgm_register/C3295  ( .a(enable), .b(a[70]), .out(
        \prgm_register/n143 ) );
  nand2 \prgm_register/C3296  ( .a(\prgm_register/en_not ), .b(a[71]), .out(
        \prgm_register/n144 ) );
  nand2 \prgm_register/C3297  ( .a(\prgm_register/n143 ), .b(
        \prgm_register/n144 ), .out(\prgm_register/or_signal [71]) );
  nand2 \prgm_register/C3298  ( .a(enable), .b(a[71]), .out(
        \prgm_register/n145 ) );
  nand2 \prgm_register/C3299  ( .a(\prgm_register/en_not ), .b(a[72]), .out(
        \prgm_register/n146 ) );
  nand2 \prgm_register/C3300  ( .a(\prgm_register/n145 ), .b(
        \prgm_register/n146 ), .out(\prgm_register/or_signal [72]) );
  nand2 \prgm_register/C3301  ( .a(enable), .b(a[72]), .out(
        \prgm_register/n147 ) );
  nand2 \prgm_register/C3302  ( .a(\prgm_register/en_not ), .b(a[73]), .out(
        \prgm_register/n148 ) );
  nand2 \prgm_register/C3303  ( .a(\prgm_register/n147 ), .b(
        \prgm_register/n148 ), .out(\prgm_register/or_signal [73]) );
  nand2 \prgm_register/C3304  ( .a(enable), .b(a[73]), .out(
        \prgm_register/n149 ) );
  nand2 \prgm_register/C3305  ( .a(\prgm_register/en_not ), .b(a[74]), .out(
        \prgm_register/n150 ) );
  nand2 \prgm_register/C3306  ( .a(\prgm_register/n149 ), .b(
        \prgm_register/n150 ), .out(\prgm_register/or_signal [74]) );
  nand2 \prgm_register/C3307  ( .a(enable), .b(a[74]), .out(
        \prgm_register/n151 ) );
  nand2 \prgm_register/C3308  ( .a(\prgm_register/en_not ), .b(a[75]), .out(
        \prgm_register/n152 ) );
  nand2 \prgm_register/C3309  ( .a(\prgm_register/n151 ), .b(
        \prgm_register/n152 ), .out(\prgm_register/or_signal [75]) );
  nand2 \prgm_register/C3310  ( .a(enable), .b(a[75]), .out(
        \prgm_register/n153 ) );
  nand2 \prgm_register/C3311  ( .a(\prgm_register/en_not ), .b(a[76]), .out(
        \prgm_register/n154 ) );
  nand2 \prgm_register/C3312  ( .a(\prgm_register/n153 ), .b(
        \prgm_register/n154 ), .out(\prgm_register/or_signal [76]) );
  nand2 \prgm_register/C3313  ( .a(enable), .b(a[76]), .out(
        \prgm_register/n155 ) );
  nand2 \prgm_register/C3314  ( .a(\prgm_register/en_not ), .b(a[77]), .out(
        \prgm_register/n156 ) );
  nand2 \prgm_register/C3315  ( .a(\prgm_register/n155 ), .b(
        \prgm_register/n156 ), .out(\prgm_register/or_signal [77]) );
  nand2 \prgm_register/C3316  ( .a(enable), .b(a[77]), .out(
        \prgm_register/n157 ) );
  nand2 \prgm_register/C3317  ( .a(\prgm_register/en_not ), .b(a[78]), .out(
        \prgm_register/n158 ) );
  nand2 \prgm_register/C3318  ( .a(\prgm_register/n157 ), .b(
        \prgm_register/n158 ), .out(\prgm_register/or_signal [78]) );
  nand2 \prgm_register/C3319  ( .a(enable), .b(a[78]), .out(
        \prgm_register/n159 ) );
  nand2 \prgm_register/C3320  ( .a(\prgm_register/en_not ), .b(a[79]), .out(
        \prgm_register/n160 ) );
  nand2 \prgm_register/C3321  ( .a(\prgm_register/n159 ), .b(
        \prgm_register/n160 ), .out(\prgm_register/or_signal [79]) );
  nand2 \prgm_register/C3322  ( .a(enable), .b(a[79]), .out(
        \prgm_register/n161 ) );
  nand2 \prgm_register/C3323  ( .a(\prgm_register/en_not ), .b(a[80]), .out(
        \prgm_register/n162 ) );
  nand2 \prgm_register/C3324  ( .a(\prgm_register/n161 ), .b(
        \prgm_register/n162 ), .out(\prgm_register/or_signal [80]) );
  nand2 \prgm_register/C3325  ( .a(enable), .b(a[80]), .out(
        \prgm_register/n163 ) );
  nand2 \prgm_register/C3326  ( .a(\prgm_register/en_not ), .b(a[81]), .out(
        \prgm_register/n164 ) );
  nand2 \prgm_register/C3327  ( .a(\prgm_register/n163 ), .b(
        \prgm_register/n164 ), .out(\prgm_register/or_signal [81]) );
  nand2 \prgm_register/C3328  ( .a(enable), .b(a[81]), .out(
        \prgm_register/n165 ) );
  nand2 \prgm_register/C3329  ( .a(\prgm_register/en_not ), .b(a[82]), .out(
        \prgm_register/n166 ) );
  nand2 \prgm_register/C3330  ( .a(\prgm_register/n165 ), .b(
        \prgm_register/n166 ), .out(\prgm_register/or_signal [82]) );
  nand2 \prgm_register/C3331  ( .a(enable), .b(a[82]), .out(
        \prgm_register/n167 ) );
  nand2 \prgm_register/C3332  ( .a(\prgm_register/en_not ), .b(a[83]), .out(
        \prgm_register/n168 ) );
  nand2 \prgm_register/C3333  ( .a(\prgm_register/n167 ), .b(
        \prgm_register/n168 ), .out(\prgm_register/or_signal [83]) );
  nand2 \prgm_register/C3334  ( .a(enable), .b(a[83]), .out(
        \prgm_register/n169 ) );
  nand2 \prgm_register/C3335  ( .a(\prgm_register/en_not ), .b(a[84]), .out(
        \prgm_register/n170 ) );
  nand2 \prgm_register/C3336  ( .a(\prgm_register/n169 ), .b(
        \prgm_register/n170 ), .out(\prgm_register/or_signal [84]) );
  nand2 \prgm_register/C3337  ( .a(enable), .b(a[84]), .out(
        \prgm_register/n171 ) );
  nand2 \prgm_register/C3338  ( .a(\prgm_register/en_not ), .b(a[85]), .out(
        \prgm_register/n172 ) );
  nand2 \prgm_register/C3339  ( .a(\prgm_register/n171 ), .b(
        \prgm_register/n172 ), .out(\prgm_register/or_signal [85]) );
  nand2 \prgm_register/C3340  ( .a(enable), .b(a[85]), .out(
        \prgm_register/n173 ) );
  nand2 \prgm_register/C3341  ( .a(\prgm_register/en_not ), .b(a[86]), .out(
        \prgm_register/n174 ) );
  nand2 \prgm_register/C3342  ( .a(\prgm_register/n173 ), .b(
        \prgm_register/n174 ), .out(\prgm_register/or_signal [86]) );
  nand2 \prgm_register/C3343  ( .a(enable), .b(a[86]), .out(
        \prgm_register/n175 ) );
  nand2 \prgm_register/C3344  ( .a(\prgm_register/en_not ), .b(a[87]), .out(
        \prgm_register/n176 ) );
  nand2 \prgm_register/C3345  ( .a(\prgm_register/n175 ), .b(
        \prgm_register/n176 ), .out(\prgm_register/or_signal [87]) );
  nand2 \prgm_register/C3346  ( .a(enable), .b(a[87]), .out(
        \prgm_register/n177 ) );
  nand2 \prgm_register/C3347  ( .a(\prgm_register/en_not ), .b(a[88]), .out(
        \prgm_register/n178 ) );
  nand2 \prgm_register/C3348  ( .a(\prgm_register/n177 ), .b(
        \prgm_register/n178 ), .out(\prgm_register/or_signal [88]) );
  nand2 \prgm_register/C3349  ( .a(enable), .b(a[88]), .out(
        \prgm_register/n179 ) );
  nand2 \prgm_register/C3350  ( .a(\prgm_register/en_not ), .b(a[89]), .out(
        \prgm_register/n180 ) );
  nand2 \prgm_register/C3351  ( .a(\prgm_register/n179 ), .b(
        \prgm_register/n180 ), .out(\prgm_register/or_signal [89]) );
  nand2 \prgm_register/C3352  ( .a(enable), .b(a[89]), .out(
        \prgm_register/n181 ) );
  nand2 \prgm_register/C3353  ( .a(\prgm_register/en_not ), .b(a[90]), .out(
        \prgm_register/n182 ) );
  nand2 \prgm_register/C3354  ( .a(\prgm_register/n181 ), .b(
        \prgm_register/n182 ), .out(\prgm_register/or_signal [90]) );
  nand2 \prgm_register/C3355  ( .a(enable), .b(a[90]), .out(
        \prgm_register/n183 ) );
  nand2 \prgm_register/C3356  ( .a(\prgm_register/en_not ), .b(a[91]), .out(
        \prgm_register/n184 ) );
  nand2 \prgm_register/C3357  ( .a(\prgm_register/n183 ), .b(
        \prgm_register/n184 ), .out(\prgm_register/or_signal [91]) );
  nand2 \prgm_register/C3358  ( .a(enable), .b(a[91]), .out(
        \prgm_register/n185 ) );
  nand2 \prgm_register/C3359  ( .a(\prgm_register/en_not ), .b(a[92]), .out(
        \prgm_register/n186 ) );
  nand2 \prgm_register/C3360  ( .a(\prgm_register/n185 ), .b(
        \prgm_register/n186 ), .out(\prgm_register/or_signal [92]) );
  nand2 \prgm_register/C3361  ( .a(enable), .b(a[92]), .out(
        \prgm_register/n187 ) );
  nand2 \prgm_register/C3362  ( .a(\prgm_register/en_not ), .b(a[93]), .out(
        \prgm_register/n188 ) );
  nand2 \prgm_register/C3363  ( .a(\prgm_register/n187 ), .b(
        \prgm_register/n188 ), .out(\prgm_register/or_signal [93]) );
  nand2 \prgm_register/C3364  ( .a(enable), .b(a[93]), .out(
        \prgm_register/n189 ) );
  nand2 \prgm_register/C3365  ( .a(\prgm_register/en_not ), .b(a[94]), .out(
        \prgm_register/n190 ) );
  nand2 \prgm_register/C3366  ( .a(\prgm_register/n189 ), .b(
        \prgm_register/n190 ), .out(\prgm_register/or_signal [94]) );
  nand2 \prgm_register/C3367  ( .a(enable), .b(a[94]), .out(
        \prgm_register/n191 ) );
  nand2 \prgm_register/C3368  ( .a(\prgm_register/en_not ), .b(a[95]), .out(
        \prgm_register/n192 ) );
  nand2 \prgm_register/C3369  ( .a(\prgm_register/n191 ), .b(
        \prgm_register/n192 ), .out(\prgm_register/or_signal [95]) );
  nand2 \prgm_register/C3370  ( .a(enable), .b(a[95]), .out(
        \prgm_register/n193 ) );
  nand2 \prgm_register/C3371  ( .a(\prgm_register/en_not ), .b(a[96]), .out(
        \prgm_register/n194 ) );
  nand2 \prgm_register/C3372  ( .a(\prgm_register/n193 ), .b(
        \prgm_register/n194 ), .out(\prgm_register/or_signal [96]) );
  nand2 \prgm_register/C3373  ( .a(enable), .b(a[96]), .out(
        \prgm_register/n195 ) );
  nand2 \prgm_register/C3374  ( .a(\prgm_register/en_not ), .b(a[97]), .out(
        \prgm_register/n196 ) );
  nand2 \prgm_register/C3375  ( .a(\prgm_register/n195 ), .b(
        \prgm_register/n196 ), .out(\prgm_register/or_signal [97]) );
  nand2 \prgm_register/C3376  ( .a(enable), .b(a[97]), .out(
        \prgm_register/n197 ) );
  nand2 \prgm_register/C3377  ( .a(\prgm_register/en_not ), .b(a[98]), .out(
        \prgm_register/n198 ) );
  nand2 \prgm_register/C3378  ( .a(\prgm_register/n197 ), .b(
        \prgm_register/n198 ), .out(\prgm_register/or_signal [98]) );
  nand2 \prgm_register/C3379  ( .a(enable), .b(a[98]), .out(
        \prgm_register/n199 ) );
  nand2 \prgm_register/C3380  ( .a(\prgm_register/en_not ), .b(a[99]), .out(
        \prgm_register/n200 ) );
  nand2 \prgm_register/C3381  ( .a(\prgm_register/n199 ), .b(
        \prgm_register/n200 ), .out(\prgm_register/or_signal [99]) );
  nand2 \prgm_register/C3382  ( .a(enable), .b(a[99]), .out(
        \prgm_register/n201 ) );
  nand2 \prgm_register/C3383  ( .a(\prgm_register/en_not ), .b(a[100]), .out(
        \prgm_register/n202 ) );
  nand2 \prgm_register/C3384  ( .a(\prgm_register/n201 ), .b(
        \prgm_register/n202 ), .out(\prgm_register/or_signal [100]) );
  nand2 \prgm_register/C3385  ( .a(enable), .b(a[100]), .out(
        \prgm_register/n203 ) );
  nand2 \prgm_register/C3386  ( .a(\prgm_register/en_not ), .b(a[101]), .out(
        \prgm_register/n204 ) );
  nand2 \prgm_register/C3387  ( .a(\prgm_register/n203 ), .b(
        \prgm_register/n204 ), .out(\prgm_register/or_signal [101]) );
  nand2 \prgm_register/C3388  ( .a(enable), .b(a[101]), .out(
        \prgm_register/n205 ) );
  nand2 \prgm_register/C3389  ( .a(\prgm_register/en_not ), .b(a[102]), .out(
        \prgm_register/n206 ) );
  nand2 \prgm_register/C3390  ( .a(\prgm_register/n205 ), .b(
        \prgm_register/n206 ), .out(\prgm_register/or_signal [102]) );
  nand2 \prgm_register/C3391  ( .a(enable), .b(a[102]), .out(
        \prgm_register/n207 ) );
  nand2 \prgm_register/C3392  ( .a(\prgm_register/en_not ), .b(a[103]), .out(
        \prgm_register/n208 ) );
  nand2 \prgm_register/C3393  ( .a(\prgm_register/n207 ), .b(
        \prgm_register/n208 ), .out(\prgm_register/or_signal [103]) );
  nand2 \prgm_register/C3394  ( .a(enable), .b(a[103]), .out(
        \prgm_register/n209 ) );
  nand2 \prgm_register/C3395  ( .a(\prgm_register/en_not ), .b(a[104]), .out(
        \prgm_register/n210 ) );
  nand2 \prgm_register/C3396  ( .a(\prgm_register/n209 ), .b(
        \prgm_register/n210 ), .out(\prgm_register/or_signal [104]) );
  nand2 \prgm_register/C3397  ( .a(enable), .b(a[104]), .out(
        \prgm_register/n211 ) );
  nand2 \prgm_register/C3398  ( .a(\prgm_register/en_not ), .b(a[105]), .out(
        \prgm_register/n212 ) );
  nand2 \prgm_register/C3399  ( .a(\prgm_register/n211 ), .b(
        \prgm_register/n212 ), .out(\prgm_register/or_signal [105]) );
  nand2 \prgm_register/C3400  ( .a(enable), .b(a[105]), .out(
        \prgm_register/n213 ) );
  nand2 \prgm_register/C3401  ( .a(\prgm_register/en_not ), .b(a[106]), .out(
        \prgm_register/n214 ) );
  nand2 \prgm_register/C3402  ( .a(\prgm_register/n213 ), .b(
        \prgm_register/n214 ), .out(\prgm_register/or_signal [106]) );
  nand2 \prgm_register/C3403  ( .a(enable), .b(a[106]), .out(
        \prgm_register/n215 ) );
  nand2 \prgm_register/C3404  ( .a(\prgm_register/en_not ), .b(a[107]), .out(
        \prgm_register/n216 ) );
  nand2 \prgm_register/C3405  ( .a(\prgm_register/n215 ), .b(
        \prgm_register/n216 ), .out(\prgm_register/or_signal [107]) );
  nand2 \prgm_register/C3406  ( .a(enable), .b(a[107]), .out(
        \prgm_register/n217 ) );
  nand2 \prgm_register/C3407  ( .a(\prgm_register/en_not ), .b(a[108]), .out(
        \prgm_register/n218 ) );
  nand2 \prgm_register/C3408  ( .a(\prgm_register/n217 ), .b(
        \prgm_register/n218 ), .out(\prgm_register/or_signal [108]) );
  nand2 \prgm_register/C3409  ( .a(enable), .b(a[108]), .out(
        \prgm_register/n219 ) );
  nand2 \prgm_register/C3410  ( .a(\prgm_register/en_not ), .b(a[109]), .out(
        \prgm_register/n220 ) );
  nand2 \prgm_register/C3411  ( .a(\prgm_register/n219 ), .b(
        \prgm_register/n220 ), .out(\prgm_register/or_signal [109]) );
  nand2 \prgm_register/C3412  ( .a(enable), .b(a[109]), .out(
        \prgm_register/n221 ) );
  nand2 \prgm_register/C3413  ( .a(\prgm_register/en_not ), .b(a[110]), .out(
        \prgm_register/n222 ) );
  nand2 \prgm_register/C3414  ( .a(\prgm_register/n221 ), .b(
        \prgm_register/n222 ), .out(\prgm_register/or_signal [110]) );
  nand2 \prgm_register/C3415  ( .a(enable), .b(a[110]), .out(
        \prgm_register/n223 ) );
  nand2 \prgm_register/C3416  ( .a(\prgm_register/en_not ), .b(a[111]), .out(
        \prgm_register/n224 ) );
  nand2 \prgm_register/C3417  ( .a(\prgm_register/n223 ), .b(
        \prgm_register/n224 ), .out(\prgm_register/or_signal [111]) );
  nand2 \prgm_register/C3418  ( .a(enable), .b(a[111]), .out(
        \prgm_register/n225 ) );
  nand2 \prgm_register/C3419  ( .a(\prgm_register/en_not ), .b(a[112]), .out(
        \prgm_register/n226 ) );
  nand2 \prgm_register/C3420  ( .a(\prgm_register/n225 ), .b(
        \prgm_register/n226 ), .out(\prgm_register/or_signal [112]) );
  nand2 \prgm_register/C3421  ( .a(enable), .b(a[112]), .out(
        \prgm_register/n227 ) );
  nand2 \prgm_register/C3422  ( .a(\prgm_register/en_not ), .b(a[113]), .out(
        \prgm_register/n228 ) );
  nand2 \prgm_register/C3423  ( .a(\prgm_register/n227 ), .b(
        \prgm_register/n228 ), .out(\prgm_register/or_signal [113]) );
  nand2 \prgm_register/C3424  ( .a(enable), .b(a[113]), .out(
        \prgm_register/n229 ) );
  nand2 \prgm_register/C3425  ( .a(\prgm_register/en_not ), .b(a[114]), .out(
        \prgm_register/n230 ) );
  nand2 \prgm_register/C3426  ( .a(\prgm_register/n229 ), .b(
        \prgm_register/n230 ), .out(\prgm_register/or_signal [114]) );
  nand2 \prgm_register/C3427  ( .a(enable), .b(a[114]), .out(
        \prgm_register/n231 ) );
  nand2 \prgm_register/C3428  ( .a(\prgm_register/en_not ), .b(a[115]), .out(
        \prgm_register/n232 ) );
  nand2 \prgm_register/C3429  ( .a(\prgm_register/n231 ), .b(
        \prgm_register/n232 ), .out(\prgm_register/or_signal [115]) );
  nand2 \prgm_register/C3430  ( .a(enable), .b(a[115]), .out(
        \prgm_register/n233 ) );
  nand2 \prgm_register/C3431  ( .a(\prgm_register/en_not ), .b(a[116]), .out(
        \prgm_register/n234 ) );
  nand2 \prgm_register/C3432  ( .a(\prgm_register/n233 ), .b(
        \prgm_register/n234 ), .out(\prgm_register/or_signal [116]) );
  nand2 \prgm_register/C3433  ( .a(enable), .b(a[116]), .out(
        \prgm_register/n235 ) );
  nand2 \prgm_register/C3434  ( .a(\prgm_register/en_not ), .b(a[117]), .out(
        \prgm_register/n236 ) );
  nand2 \prgm_register/C3435  ( .a(\prgm_register/n235 ), .b(
        \prgm_register/n236 ), .out(\prgm_register/or_signal [117]) );
  nand2 \prgm_register/C3436  ( .a(enable), .b(a[117]), .out(
        \prgm_register/n237 ) );
  nand2 \prgm_register/C3437  ( .a(\prgm_register/en_not ), .b(a[118]), .out(
        \prgm_register/n238 ) );
  nand2 \prgm_register/C3438  ( .a(\prgm_register/n237 ), .b(
        \prgm_register/n238 ), .out(\prgm_register/or_signal [118]) );
  nand2 \prgm_register/C3439  ( .a(enable), .b(a[118]), .out(
        \prgm_register/n239 ) );
  nand2 \prgm_register/C3440  ( .a(\prgm_register/en_not ), .b(a[119]), .out(
        \prgm_register/n240 ) );
  nand2 \prgm_register/C3441  ( .a(\prgm_register/n239 ), .b(
        \prgm_register/n240 ), .out(\prgm_register/or_signal [119]) );
  nand2 \prgm_register/C3442  ( .a(enable), .b(a[119]), .out(
        \prgm_register/n241 ) );
  nand2 \prgm_register/C3443  ( .a(\prgm_register/en_not ), .b(a[120]), .out(
        \prgm_register/n242 ) );
  nand2 \prgm_register/C3444  ( .a(\prgm_register/n241 ), .b(
        \prgm_register/n242 ), .out(\prgm_register/or_signal [120]) );
  nand2 \prgm_register/C3445  ( .a(enable), .b(a[120]), .out(
        \prgm_register/n243 ) );
  nand2 \prgm_register/C3446  ( .a(\prgm_register/en_not ), .b(a[121]), .out(
        \prgm_register/n244 ) );
  nand2 \prgm_register/C3447  ( .a(\prgm_register/n243 ), .b(
        \prgm_register/n244 ), .out(\prgm_register/or_signal [121]) );
  nand2 \prgm_register/C3448  ( .a(enable), .b(a[121]), .out(
        \prgm_register/n245 ) );
  nand2 \prgm_register/C3449  ( .a(\prgm_register/en_not ), .b(a[122]), .out(
        \prgm_register/n246 ) );
  nand2 \prgm_register/C3450  ( .a(\prgm_register/n245 ), .b(
        \prgm_register/n246 ), .out(\prgm_register/or_signal [122]) );
  nand2 \prgm_register/C3451  ( .a(enable), .b(a[122]), .out(
        \prgm_register/n247 ) );
  nand2 \prgm_register/C3452  ( .a(\prgm_register/en_not ), .b(a[123]), .out(
        \prgm_register/n248 ) );
  nand2 \prgm_register/C3453  ( .a(\prgm_register/n247 ), .b(
        \prgm_register/n248 ), .out(\prgm_register/or_signal [123]) );
  nand2 \prgm_register/C3454  ( .a(enable), .b(a[123]), .out(
        \prgm_register/n249 ) );
  nand2 \prgm_register/C3455  ( .a(\prgm_register/en_not ), .b(a[124]), .out(
        \prgm_register/n250 ) );
  nand2 \prgm_register/C3456  ( .a(\prgm_register/n249 ), .b(
        \prgm_register/n250 ), .out(\prgm_register/or_signal [124]) );
  nand2 \prgm_register/C3457  ( .a(enable), .b(a[124]), .out(
        \prgm_register/n251 ) );
  nand2 \prgm_register/C3458  ( .a(\prgm_register/en_not ), .b(a[125]), .out(
        \prgm_register/n252 ) );
  nand2 \prgm_register/C3459  ( .a(\prgm_register/n251 ), .b(
        \prgm_register/n252 ), .out(\prgm_register/or_signal [125]) );
  nand2 \prgm_register/C3460  ( .a(enable), .b(a[125]), .out(
        \prgm_register/n253 ) );
  nand2 \prgm_register/C3461  ( .a(\prgm_register/en_not ), .b(a[126]), .out(
        \prgm_register/n254 ) );
  nand2 \prgm_register/C3462  ( .a(\prgm_register/n253 ), .b(
        \prgm_register/n254 ), .out(\prgm_register/or_signal [126]) );
  nand2 \prgm_register/C3463  ( .a(enable), .b(a[126]), .out(
        \prgm_register/n255 ) );
  nand2 \prgm_register/C3464  ( .a(\prgm_register/en_not ), .b(a[127]), .out(
        \prgm_register/n256 ) );
  nand2 \prgm_register/C3465  ( .a(\prgm_register/n255 ), .b(
        \prgm_register/n256 ), .out(\prgm_register/or_signal [127]) );
  nand2 \prgm_register/C3466  ( .a(enable), .b(a[127]), .out(
        \prgm_register/n257 ) );
  nand2 \prgm_register/C3467  ( .a(\prgm_register/en_not ), .b(a[128]), .out(
        \prgm_register/n258 ) );
  nand2 \prgm_register/C3468  ( .a(\prgm_register/n257 ), .b(
        \prgm_register/n258 ), .out(\prgm_register/or_signal [128]) );
  nand2 \prgm_register/C3469  ( .a(enable), .b(a[128]), .out(
        \prgm_register/n259 ) );
  nand2 \prgm_register/C3470  ( .a(\prgm_register/en_not ), .b(a[129]), .out(
        \prgm_register/n260 ) );
  nand2 \prgm_register/C3471  ( .a(\prgm_register/n259 ), .b(
        \prgm_register/n260 ), .out(\prgm_register/or_signal [129]) );
  nand2 \prgm_register/C3472  ( .a(enable), .b(a[129]), .out(
        \prgm_register/n261 ) );
  nand2 \prgm_register/C3473  ( .a(\prgm_register/en_not ), .b(a[130]), .out(
        \prgm_register/n262 ) );
  nand2 \prgm_register/C3474  ( .a(\prgm_register/n261 ), .b(
        \prgm_register/n262 ), .out(\prgm_register/or_signal [130]) );
  nand2 \prgm_register/C3475  ( .a(enable), .b(a[130]), .out(
        \prgm_register/n263 ) );
  nand2 \prgm_register/C3476  ( .a(\prgm_register/en_not ), .b(a[131]), .out(
        \prgm_register/n264 ) );
  nand2 \prgm_register/C3477  ( .a(\prgm_register/n263 ), .b(
        \prgm_register/n264 ), .out(\prgm_register/or_signal [131]) );
  nand2 \prgm_register/C3478  ( .a(enable), .b(a[131]), .out(
        \prgm_register/n265 ) );
  nand2 \prgm_register/C3479  ( .a(\prgm_register/en_not ), .b(a[132]), .out(
        \prgm_register/n266 ) );
  nand2 \prgm_register/C3480  ( .a(\prgm_register/n265 ), .b(
        \prgm_register/n266 ), .out(\prgm_register/or_signal [132]) );
  nand2 \prgm_register/C3481  ( .a(enable), .b(a[132]), .out(
        \prgm_register/n267 ) );
  nand2 \prgm_register/C3482  ( .a(\prgm_register/en_not ), .b(a[133]), .out(
        \prgm_register/n268 ) );
  nand2 \prgm_register/C3483  ( .a(\prgm_register/n267 ), .b(
        \prgm_register/n268 ), .out(\prgm_register/or_signal [133]) );
  nand2 \prgm_register/C3484  ( .a(enable), .b(a[133]), .out(
        \prgm_register/n269 ) );
  nand2 \prgm_register/C3485  ( .a(\prgm_register/en_not ), .b(a[134]), .out(
        \prgm_register/n270 ) );
  nand2 \prgm_register/C3486  ( .a(\prgm_register/n269 ), .b(
        \prgm_register/n270 ), .out(\prgm_register/or_signal [134]) );
  nand2 \prgm_register/C3487  ( .a(enable), .b(a[134]), .out(
        \prgm_register/n271 ) );
  nand2 \prgm_register/C3488  ( .a(\prgm_register/en_not ), .b(a[135]), .out(
        \prgm_register/n272 ) );
  nand2 \prgm_register/C3489  ( .a(\prgm_register/n271 ), .b(
        \prgm_register/n272 ), .out(\prgm_register/or_signal [135]) );
  nand2 \prgm_register/C3490  ( .a(enable), .b(a[135]), .out(
        \prgm_register/n273 ) );
  nand2 \prgm_register/C3491  ( .a(\prgm_register/en_not ), .b(a[136]), .out(
        \prgm_register/n274 ) );
  nand2 \prgm_register/C3492  ( .a(\prgm_register/n273 ), .b(
        \prgm_register/n274 ), .out(\prgm_register/or_signal [136]) );
  nand2 \prgm_register/C3493  ( .a(enable), .b(a[136]), .out(
        \prgm_register/n275 ) );
  nand2 \prgm_register/C3494  ( .a(\prgm_register/en_not ), .b(a[137]), .out(
        \prgm_register/n276 ) );
  nand2 \prgm_register/C3495  ( .a(\prgm_register/n275 ), .b(
        \prgm_register/n276 ), .out(\prgm_register/or_signal [137]) );
  nand2 \prgm_register/C3496  ( .a(enable), .b(a[137]), .out(
        \prgm_register/n277 ) );
  nand2 \prgm_register/C3497  ( .a(\prgm_register/en_not ), .b(a[138]), .out(
        \prgm_register/n278 ) );
  nand2 \prgm_register/C3498  ( .a(\prgm_register/n277 ), .b(
        \prgm_register/n278 ), .out(\prgm_register/or_signal [138]) );
  nand2 \prgm_register/C3499  ( .a(enable), .b(a[138]), .out(
        \prgm_register/n279 ) );
  nand2 \prgm_register/C3500  ( .a(\prgm_register/en_not ), .b(a[139]), .out(
        \prgm_register/n280 ) );
  nand2 \prgm_register/C3501  ( .a(\prgm_register/n279 ), .b(
        \prgm_register/n280 ), .out(\prgm_register/or_signal [139]) );
  nand2 \prgm_register/C3502  ( .a(enable), .b(a[139]), .out(
        \prgm_register/n281 ) );
  nand2 \prgm_register/C3503  ( .a(\prgm_register/en_not ), .b(a[140]), .out(
        \prgm_register/n282 ) );
  nand2 \prgm_register/C3504  ( .a(\prgm_register/n281 ), .b(
        \prgm_register/n282 ), .out(\prgm_register/or_signal [140]) );
  nand2 \prgm_register/C3505  ( .a(enable), .b(a[140]), .out(
        \prgm_register/n283 ) );
  nand2 \prgm_register/C3506  ( .a(\prgm_register/en_not ), .b(a[141]), .out(
        \prgm_register/n284 ) );
  nand2 \prgm_register/C3507  ( .a(\prgm_register/n283 ), .b(
        \prgm_register/n284 ), .out(\prgm_register/or_signal [141]) );
  nand2 \prgm_register/C3508  ( .a(enable), .b(a[141]), .out(
        \prgm_register/n285 ) );
  nand2 \prgm_register/C3509  ( .a(\prgm_register/en_not ), .b(a[142]), .out(
        \prgm_register/n286 ) );
  nand2 \prgm_register/C3510  ( .a(\prgm_register/n285 ), .b(
        \prgm_register/n286 ), .out(\prgm_register/or_signal [142]) );
  nand2 \prgm_register/C3511  ( .a(enable), .b(a[142]), .out(
        \prgm_register/n287 ) );
  nand2 \prgm_register/C3512  ( .a(\prgm_register/en_not ), .b(a[143]), .out(
        \prgm_register/n288 ) );
  nand2 \prgm_register/C3513  ( .a(\prgm_register/n287 ), .b(
        \prgm_register/n288 ), .out(\prgm_register/or_signal [143]) );
  nand2 \prgm_register/C3514  ( .a(enable), .b(a[143]), .out(
        \prgm_register/n289 ) );
  nand2 \prgm_register/C3515  ( .a(\prgm_register/en_not ), .b(a[144]), .out(
        \prgm_register/n290 ) );
  nand2 \prgm_register/C3516  ( .a(\prgm_register/n289 ), .b(
        \prgm_register/n290 ), .out(\prgm_register/or_signal [144]) );
  nand2 \prgm_register/C3517  ( .a(enable), .b(a[144]), .out(
        \prgm_register/n291 ) );
  nand2 \prgm_register/C3518  ( .a(\prgm_register/en_not ), .b(a[145]), .out(
        \prgm_register/n292 ) );
  nand2 \prgm_register/C3519  ( .a(\prgm_register/n291 ), .b(
        \prgm_register/n292 ), .out(\prgm_register/or_signal [145]) );
  nand2 \prgm_register/C3520  ( .a(enable), .b(a[145]), .out(
        \prgm_register/n293 ) );
  nand2 \prgm_register/C3521  ( .a(\prgm_register/en_not ), .b(a[146]), .out(
        \prgm_register/n294 ) );
  nand2 \prgm_register/C3522  ( .a(\prgm_register/n293 ), .b(
        \prgm_register/n294 ), .out(\prgm_register/or_signal [146]) );
  nand2 \prgm_register/C3523  ( .a(enable), .b(a[146]), .out(
        \prgm_register/n295 ) );
  nand2 \prgm_register/C3524  ( .a(\prgm_register/en_not ), .b(a[147]), .out(
        \prgm_register/n296 ) );
  nand2 \prgm_register/C3525  ( .a(\prgm_register/n295 ), .b(
        \prgm_register/n296 ), .out(\prgm_register/or_signal [147]) );
  nand2 \prgm_register/C3526  ( .a(enable), .b(a[147]), .out(
        \prgm_register/n297 ) );
  nand2 \prgm_register/C3527  ( .a(\prgm_register/en_not ), .b(a[148]), .out(
        \prgm_register/n298 ) );
  nand2 \prgm_register/C3528  ( .a(\prgm_register/n297 ), .b(
        \prgm_register/n298 ), .out(\prgm_register/or_signal [148]) );
  nand2 \prgm_register/C3529  ( .a(enable), .b(a[148]), .out(
        \prgm_register/n299 ) );
  nand2 \prgm_register/C3530  ( .a(\prgm_register/en_not ), .b(a[149]), .out(
        \prgm_register/n300 ) );
  nand2 \prgm_register/C3531  ( .a(\prgm_register/n299 ), .b(
        \prgm_register/n300 ), .out(\prgm_register/or_signal [149]) );
  nand2 \prgm_register/C3532  ( .a(enable), .b(a[149]), .out(
        \prgm_register/n301 ) );
  nand2 \prgm_register/C3533  ( .a(\prgm_register/en_not ), .b(a[150]), .out(
        \prgm_register/n302 ) );
  nand2 \prgm_register/C3534  ( .a(\prgm_register/n301 ), .b(
        \prgm_register/n302 ), .out(\prgm_register/or_signal [150]) );
  nand2 \prgm_register/C3535  ( .a(enable), .b(a[150]), .out(
        \prgm_register/n303 ) );
  nand2 \prgm_register/C3536  ( .a(\prgm_register/en_not ), .b(a[151]), .out(
        \prgm_register/n304 ) );
  nand2 \prgm_register/C3537  ( .a(\prgm_register/n303 ), .b(
        \prgm_register/n304 ), .out(\prgm_register/or_signal [151]) );
  nand2 \prgm_register/C3538  ( .a(enable), .b(a[151]), .out(
        \prgm_register/n305 ) );
  nand2 \prgm_register/C3539  ( .a(\prgm_register/en_not ), .b(a[152]), .out(
        \prgm_register/n306 ) );
  nand2 \prgm_register/C3540  ( .a(\prgm_register/n305 ), .b(
        \prgm_register/n306 ), .out(\prgm_register/or_signal [152]) );
  nand2 \prgm_register/C3541  ( .a(enable), .b(a[152]), .out(
        \prgm_register/n307 ) );
  nand2 \prgm_register/C3542  ( .a(\prgm_register/en_not ), .b(a[153]), .out(
        \prgm_register/n308 ) );
  nand2 \prgm_register/C3543  ( .a(\prgm_register/n307 ), .b(
        \prgm_register/n308 ), .out(\prgm_register/or_signal [153]) );
  nand2 \prgm_register/C3544  ( .a(enable), .b(a[153]), .out(
        \prgm_register/n309 ) );
  nand2 \prgm_register/C3545  ( .a(\prgm_register/en_not ), .b(a[154]), .out(
        \prgm_register/n310 ) );
  nand2 \prgm_register/C3546  ( .a(\prgm_register/n309 ), .b(
        \prgm_register/n310 ), .out(\prgm_register/or_signal [154]) );
  nand2 \prgm_register/C3547  ( .a(enable), .b(a[154]), .out(
        \prgm_register/n311 ) );
  nand2 \prgm_register/C3548  ( .a(\prgm_register/en_not ), .b(a[155]), .out(
        \prgm_register/n312 ) );
  nand2 \prgm_register/C3549  ( .a(\prgm_register/n311 ), .b(
        \prgm_register/n312 ), .out(\prgm_register/or_signal [155]) );
  nand2 \prgm_register/C3550  ( .a(enable), .b(a[155]), .out(
        \prgm_register/n313 ) );
  nand2 \prgm_register/C3551  ( .a(\prgm_register/en_not ), .b(a[156]), .out(
        \prgm_register/n314 ) );
  nand2 \prgm_register/C3552  ( .a(\prgm_register/n313 ), .b(
        \prgm_register/n314 ), .out(\prgm_register/or_signal [156]) );
  nand2 \prgm_register/C3553  ( .a(enable), .b(a[156]), .out(
        \prgm_register/n315 ) );
  nand2 \prgm_register/C3554  ( .a(\prgm_register/en_not ), .b(a[157]), .out(
        \prgm_register/n316 ) );
  nand2 \prgm_register/C3555  ( .a(\prgm_register/n315 ), .b(
        \prgm_register/n316 ), .out(\prgm_register/or_signal [157]) );
  nand2 \prgm_register/C3556  ( .a(enable), .b(a[157]), .out(
        \prgm_register/n317 ) );
  nand2 \prgm_register/C3557  ( .a(\prgm_register/en_not ), .b(a[158]), .out(
        \prgm_register/n318 ) );
  nand2 \prgm_register/C3558  ( .a(\prgm_register/n317 ), .b(
        \prgm_register/n318 ), .out(\prgm_register/or_signal [158]) );
  nand2 \prgm_register/C3559  ( .a(enable), .b(a[158]), .out(
        \prgm_register/n319 ) );
  nand2 \prgm_register/C3560  ( .a(\prgm_register/en_not ), .b(a[159]), .out(
        \prgm_register/n320 ) );
  nand2 \prgm_register/C3561  ( .a(\prgm_register/n319 ), .b(
        \prgm_register/n320 ), .out(\prgm_register/or_signal [159]) );
  nand2 \prgm_register/C3562  ( .a(enable), .b(a[159]), .out(
        \prgm_register/n321 ) );
  nand2 \prgm_register/C3563  ( .a(\prgm_register/en_not ), .b(a[160]), .out(
        \prgm_register/n322 ) );
  nand2 \prgm_register/C3564  ( .a(\prgm_register/n321 ), .b(
        \prgm_register/n322 ), .out(\prgm_register/or_signal [160]) );
  nand2 \prgm_register/C3565  ( .a(enable), .b(a[160]), .out(
        \prgm_register/n323 ) );
  nand2 \prgm_register/C3566  ( .a(\prgm_register/en_not ), .b(a[161]), .out(
        \prgm_register/n324 ) );
  nand2 \prgm_register/C3567  ( .a(\prgm_register/n323 ), .b(
        \prgm_register/n324 ), .out(\prgm_register/or_signal [161]) );
  nand2 \prgm_register/C3568  ( .a(enable), .b(a[161]), .out(
        \prgm_register/n325 ) );
  nand2 \prgm_register/C3569  ( .a(\prgm_register/en_not ), .b(a[162]), .out(
        \prgm_register/n326 ) );
  nand2 \prgm_register/C3570  ( .a(\prgm_register/n325 ), .b(
        \prgm_register/n326 ), .out(\prgm_register/or_signal [162]) );
  nand2 \prgm_register/C3571  ( .a(enable), .b(a[162]), .out(
        \prgm_register/n327 ) );
  nand2 \prgm_register/C3572  ( .a(\prgm_register/en_not ), .b(a[163]), .out(
        \prgm_register/n328 ) );
  nand2 \prgm_register/C3573  ( .a(\prgm_register/n327 ), .b(
        \prgm_register/n328 ), .out(\prgm_register/or_signal [163]) );
  nand2 \prgm_register/C3574  ( .a(enable), .b(a[163]), .out(
        \prgm_register/n329 ) );
  nand2 \prgm_register/C3575  ( .a(\prgm_register/en_not ), .b(a[164]), .out(
        \prgm_register/n330 ) );
  nand2 \prgm_register/C3576  ( .a(\prgm_register/n329 ), .b(
        \prgm_register/n330 ), .out(\prgm_register/or_signal [164]) );
  nand2 \prgm_register/C3577  ( .a(enable), .b(a[164]), .out(
        \prgm_register/n331 ) );
  nand2 \prgm_register/C3578  ( .a(\prgm_register/en_not ), .b(a[165]), .out(
        \prgm_register/n332 ) );
  nand2 \prgm_register/C3579  ( .a(\prgm_register/n331 ), .b(
        \prgm_register/n332 ), .out(\prgm_register/or_signal [165]) );
  nand2 \prgm_register/C3580  ( .a(enable), .b(a[165]), .out(
        \prgm_register/n333 ) );
  nand2 \prgm_register/C3581  ( .a(\prgm_register/en_not ), .b(a[166]), .out(
        \prgm_register/n334 ) );
  nand2 \prgm_register/C3582  ( .a(\prgm_register/n333 ), .b(
        \prgm_register/n334 ), .out(\prgm_register/or_signal [166]) );
  nand2 \prgm_register/C3583  ( .a(enable), .b(a[166]), .out(
        \prgm_register/n335 ) );
  nand2 \prgm_register/C3584  ( .a(\prgm_register/en_not ), .b(a[167]), .out(
        \prgm_register/n336 ) );
  nand2 \prgm_register/C3585  ( .a(\prgm_register/n335 ), .b(
        \prgm_register/n336 ), .out(\prgm_register/or_signal [167]) );
  nand2 \prgm_register/C3586  ( .a(enable), .b(a[167]), .out(
        \prgm_register/n337 ) );
  nand2 \prgm_register/C3587  ( .a(\prgm_register/en_not ), .b(a[168]), .out(
        \prgm_register/n338 ) );
  nand2 \prgm_register/C3588  ( .a(\prgm_register/n337 ), .b(
        \prgm_register/n338 ), .out(\prgm_register/or_signal [168]) );
  nand2 \prgm_register/C3589  ( .a(enable), .b(a[168]), .out(
        \prgm_register/n339 ) );
  nand2 \prgm_register/C3590  ( .a(\prgm_register/en_not ), .b(a[169]), .out(
        \prgm_register/n340 ) );
  nand2 \prgm_register/C3591  ( .a(\prgm_register/n339 ), .b(
        \prgm_register/n340 ), .out(\prgm_register/or_signal [169]) );
  nand2 \prgm_register/C3592  ( .a(enable), .b(a[169]), .out(
        \prgm_register/n341 ) );
  nand2 \prgm_register/C3593  ( .a(\prgm_register/en_not ), .b(a[170]), .out(
        \prgm_register/n342 ) );
  nand2 \prgm_register/C3594  ( .a(\prgm_register/n341 ), .b(
        \prgm_register/n342 ), .out(\prgm_register/or_signal [170]) );
  nand2 \prgm_register/C3595  ( .a(enable), .b(a[170]), .out(
        \prgm_register/n343 ) );
  nand2 \prgm_register/C3596  ( .a(\prgm_register/en_not ), .b(a[171]), .out(
        \prgm_register/n344 ) );
  nand2 \prgm_register/C3597  ( .a(\prgm_register/n343 ), .b(
        \prgm_register/n344 ), .out(\prgm_register/or_signal [171]) );
  nand2 \prgm_register/C3598  ( .a(enable), .b(a[171]), .out(
        \prgm_register/n345 ) );
  nand2 \prgm_register/C3599  ( .a(\prgm_register/en_not ), .b(a[172]), .out(
        \prgm_register/n346 ) );
  nand2 \prgm_register/C3600  ( .a(\prgm_register/n345 ), .b(
        \prgm_register/n346 ), .out(\prgm_register/or_signal [172]) );
  nand2 \prgm_register/C3601  ( .a(enable), .b(a[172]), .out(
        \prgm_register/n347 ) );
  nand2 \prgm_register/C3602  ( .a(\prgm_register/en_not ), .b(a[173]), .out(
        \prgm_register/n348 ) );
  nand2 \prgm_register/C3603  ( .a(\prgm_register/n347 ), .b(
        \prgm_register/n348 ), .out(\prgm_register/or_signal [173]) );
  nand2 \prgm_register/C3604  ( .a(enable), .b(a[173]), .out(
        \prgm_register/n349 ) );
  nand2 \prgm_register/C3605  ( .a(\prgm_register/en_not ), .b(a[174]), .out(
        \prgm_register/n350 ) );
  nand2 \prgm_register/C3606  ( .a(\prgm_register/n349 ), .b(
        \prgm_register/n350 ), .out(\prgm_register/or_signal [174]) );
  nand2 \prgm_register/C3607  ( .a(enable), .b(a[174]), .out(
        \prgm_register/n351 ) );
  nand2 \prgm_register/C3608  ( .a(\prgm_register/en_not ), .b(a[175]), .out(
        \prgm_register/n352 ) );
  nand2 \prgm_register/C3609  ( .a(\prgm_register/n351 ), .b(
        \prgm_register/n352 ), .out(\prgm_register/or_signal [175]) );
  nand2 \prgm_register/C3610  ( .a(enable), .b(a[175]), .out(
        \prgm_register/n353 ) );
  nand2 \prgm_register/C3611  ( .a(\prgm_register/en_not ), .b(a[176]), .out(
        \prgm_register/n354 ) );
  nand2 \prgm_register/C3612  ( .a(\prgm_register/n353 ), .b(
        \prgm_register/n354 ), .out(\prgm_register/or_signal [176]) );
  nand2 \prgm_register/C3613  ( .a(enable), .b(a[176]), .out(
        \prgm_register/n355 ) );
  nand2 \prgm_register/C3614  ( .a(\prgm_register/en_not ), .b(a[177]), .out(
        \prgm_register/n356 ) );
  nand2 \prgm_register/C3615  ( .a(\prgm_register/n355 ), .b(
        \prgm_register/n356 ), .out(\prgm_register/or_signal [177]) );
  nand2 \prgm_register/C3616  ( .a(enable), .b(a[177]), .out(
        \prgm_register/n357 ) );
  nand2 \prgm_register/C3617  ( .a(\prgm_register/en_not ), .b(a[178]), .out(
        \prgm_register/n358 ) );
  nand2 \prgm_register/C3618  ( .a(\prgm_register/n357 ), .b(
        \prgm_register/n358 ), .out(\prgm_register/or_signal [178]) );
  nand2 \prgm_register/C3619  ( .a(enable), .b(a[178]), .out(
        \prgm_register/n359 ) );
  nand2 \prgm_register/C3620  ( .a(\prgm_register/en_not ), .b(a[179]), .out(
        \prgm_register/n360 ) );
  nand2 \prgm_register/C3621  ( .a(\prgm_register/n359 ), .b(
        \prgm_register/n360 ), .out(\prgm_register/or_signal [179]) );
  nand2 \prgm_register/C3622  ( .a(enable), .b(a[179]), .out(
        \prgm_register/n361 ) );
  nand2 \prgm_register/C3623  ( .a(\prgm_register/en_not ), .b(a[180]), .out(
        \prgm_register/n362 ) );
  nand2 \prgm_register/C3624  ( .a(\prgm_register/n361 ), .b(
        \prgm_register/n362 ), .out(\prgm_register/or_signal [180]) );
  nand2 \prgm_register/C3625  ( .a(enable), .b(a[180]), .out(
        \prgm_register/n363 ) );
  nand2 \prgm_register/C3626  ( .a(\prgm_register/en_not ), .b(a[181]), .out(
        \prgm_register/n364 ) );
  nand2 \prgm_register/C3627  ( .a(\prgm_register/n363 ), .b(
        \prgm_register/n364 ), .out(\prgm_register/or_signal [181]) );
  nand2 \prgm_register/C3628  ( .a(enable), .b(a[181]), .out(
        \prgm_register/n365 ) );
  nand2 \prgm_register/C3629  ( .a(\prgm_register/en_not ), .b(a[182]), .out(
        \prgm_register/n366 ) );
  nand2 \prgm_register/C3630  ( .a(\prgm_register/n365 ), .b(
        \prgm_register/n366 ), .out(\prgm_register/or_signal [182]) );
  nand2 \prgm_register/C3631  ( .a(enable), .b(a[182]), .out(
        \prgm_register/n367 ) );
  nand2 \prgm_register/C3632  ( .a(\prgm_register/en_not ), .b(a[183]), .out(
        \prgm_register/n368 ) );
  nand2 \prgm_register/C3633  ( .a(\prgm_register/n367 ), .b(
        \prgm_register/n368 ), .out(\prgm_register/or_signal [183]) );
  nand2 \prgm_register/C3634  ( .a(enable), .b(a[183]), .out(
        \prgm_register/n369 ) );
  nand2 \prgm_register/C3635  ( .a(\prgm_register/en_not ), .b(a[184]), .out(
        \prgm_register/n370 ) );
  nand2 \prgm_register/C3636  ( .a(\prgm_register/n369 ), .b(
        \prgm_register/n370 ), .out(\prgm_register/or_signal [184]) );
  nand2 \prgm_register/C3637  ( .a(enable), .b(a[184]), .out(
        \prgm_register/n371 ) );
  nand2 \prgm_register/C3638  ( .a(\prgm_register/en_not ), .b(a[185]), .out(
        \prgm_register/n372 ) );
  nand2 \prgm_register/C3639  ( .a(\prgm_register/n371 ), .b(
        \prgm_register/n372 ), .out(\prgm_register/or_signal [185]) );
  nand2 \prgm_register/C3640  ( .a(enable), .b(a[185]), .out(
        \prgm_register/n373 ) );
  nand2 \prgm_register/C3641  ( .a(\prgm_register/en_not ), .b(a[186]), .out(
        \prgm_register/n374 ) );
  nand2 \prgm_register/C3642  ( .a(\prgm_register/n373 ), .b(
        \prgm_register/n374 ), .out(\prgm_register/or_signal [186]) );
  nand2 \prgm_register/C3643  ( .a(enable), .b(a[186]), .out(
        \prgm_register/n375 ) );
  nand2 \prgm_register/C3644  ( .a(\prgm_register/en_not ), .b(a[187]), .out(
        \prgm_register/n376 ) );
  nand2 \prgm_register/C3645  ( .a(\prgm_register/n375 ), .b(
        \prgm_register/n376 ), .out(\prgm_register/or_signal [187]) );
  nand2 \prgm_register/C3646  ( .a(enable), .b(a[187]), .out(
        \prgm_register/n377 ) );
  nand2 \prgm_register/C3647  ( .a(\prgm_register/en_not ), .b(a[188]), .out(
        \prgm_register/n378 ) );
  nand2 \prgm_register/C3648  ( .a(\prgm_register/n377 ), .b(
        \prgm_register/n378 ), .out(\prgm_register/or_signal [188]) );
  nand2 \prgm_register/C3649  ( .a(enable), .b(a[188]), .out(
        \prgm_register/n379 ) );
  nand2 \prgm_register/C3650  ( .a(\prgm_register/en_not ), .b(a[189]), .out(
        \prgm_register/n380 ) );
  nand2 \prgm_register/C3651  ( .a(\prgm_register/n379 ), .b(
        \prgm_register/n380 ), .out(\prgm_register/or_signal [189]) );
  nand2 \prgm_register/C3652  ( .a(enable), .b(a[189]), .out(
        \prgm_register/n381 ) );
  nand2 \prgm_register/C3653  ( .a(\prgm_register/en_not ), .b(a[190]), .out(
        \prgm_register/n382 ) );
  nand2 \prgm_register/C3654  ( .a(\prgm_register/n381 ), .b(
        \prgm_register/n382 ), .out(\prgm_register/or_signal [190]) );
  nand2 \prgm_register/C3655  ( .a(enable), .b(a[190]), .out(
        \prgm_register/n383 ) );
  nand2 \prgm_register/C3656  ( .a(\prgm_register/en_not ), .b(a[191]), .out(
        \prgm_register/n384 ) );
  nand2 \prgm_register/C3657  ( .a(\prgm_register/n383 ), .b(
        \prgm_register/n384 ), .out(\prgm_register/or_signal [191]) );
  nand2 \prgm_register/C3658  ( .a(enable), .b(a[191]), .out(
        \prgm_register/n385 ) );
  nand2 \prgm_register/C3659  ( .a(\prgm_register/en_not ), .b(a[192]), .out(
        \prgm_register/n386 ) );
  nand2 \prgm_register/C3660  ( .a(\prgm_register/n385 ), .b(
        \prgm_register/n386 ), .out(\prgm_register/or_signal [192]) );
  nand2 \prgm_register/C3661  ( .a(enable), .b(a[192]), .out(
        \prgm_register/n387 ) );
  nand2 \prgm_register/C3662  ( .a(\prgm_register/en_not ), .b(a[193]), .out(
        \prgm_register/n388 ) );
  nand2 \prgm_register/C3663  ( .a(\prgm_register/n387 ), .b(
        \prgm_register/n388 ), .out(\prgm_register/or_signal [193]) );
  nand2 \prgm_register/C3664  ( .a(enable), .b(a[193]), .out(
        \prgm_register/n389 ) );
  nand2 \prgm_register/C3665  ( .a(\prgm_register/en_not ), .b(a[194]), .out(
        \prgm_register/n390 ) );
  nand2 \prgm_register/C3666  ( .a(\prgm_register/n389 ), .b(
        \prgm_register/n390 ), .out(\prgm_register/or_signal [194]) );
  nand2 \prgm_register/C3667  ( .a(enable), .b(a[194]), .out(
        \prgm_register/n391 ) );
  nand2 \prgm_register/C3668  ( .a(\prgm_register/en_not ), .b(a[195]), .out(
        \prgm_register/n392 ) );
  nand2 \prgm_register/C3669  ( .a(\prgm_register/n391 ), .b(
        \prgm_register/n392 ), .out(\prgm_register/or_signal [195]) );
  nand2 \prgm_register/C3670  ( .a(enable), .b(a[195]), .out(
        \prgm_register/n393 ) );
  nand2 \prgm_register/C3671  ( .a(\prgm_register/en_not ), .b(a[196]), .out(
        \prgm_register/n394 ) );
  nand2 \prgm_register/C3672  ( .a(\prgm_register/n393 ), .b(
        \prgm_register/n394 ), .out(\prgm_register/or_signal [196]) );
  nand2 \prgm_register/C3673  ( .a(enable), .b(a[196]), .out(
        \prgm_register/n395 ) );
  nand2 \prgm_register/C3674  ( .a(\prgm_register/en_not ), .b(a[197]), .out(
        \prgm_register/n396 ) );
  nand2 \prgm_register/C3675  ( .a(\prgm_register/n395 ), .b(
        \prgm_register/n396 ), .out(\prgm_register/or_signal [197]) );
  nand2 \prgm_register/C3676  ( .a(enable), .b(a[197]), .out(
        \prgm_register/n397 ) );
  nand2 \prgm_register/C3677  ( .a(\prgm_register/en_not ), .b(a[198]), .out(
        \prgm_register/n398 ) );
  nand2 \prgm_register/C3678  ( .a(\prgm_register/n397 ), .b(
        \prgm_register/n398 ), .out(\prgm_register/or_signal [198]) );
  nand2 \prgm_register/C3679  ( .a(enable), .b(a[198]), .out(
        \prgm_register/n399 ) );
  nand2 \prgm_register/C3680  ( .a(\prgm_register/en_not ), .b(a[199]), .out(
        \prgm_register/n400 ) );
  nand2 \prgm_register/C3681  ( .a(\prgm_register/n399 ), .b(
        \prgm_register/n400 ), .out(\prgm_register/or_signal [199]) );
  nand2 \prgm_register/C3682  ( .a(enable), .b(a[199]), .out(
        \prgm_register/n401 ) );
  nand2 \prgm_register/C3683  ( .a(\prgm_register/en_not ), .b(a[200]), .out(
        \prgm_register/n402 ) );
  nand2 \prgm_register/C3684  ( .a(\prgm_register/n401 ), .b(
        \prgm_register/n402 ), .out(\prgm_register/or_signal [200]) );
  nand2 \prgm_register/C3685  ( .a(enable), .b(a[200]), .out(
        \prgm_register/n403 ) );
  nand2 \prgm_register/C3686  ( .a(\prgm_register/en_not ), .b(a[201]), .out(
        \prgm_register/n404 ) );
  nand2 \prgm_register/C3687  ( .a(\prgm_register/n403 ), .b(
        \prgm_register/n404 ), .out(\prgm_register/or_signal [201]) );
  nand2 \prgm_register/C3688  ( .a(enable), .b(a[201]), .out(
        \prgm_register/n405 ) );
  nand2 \prgm_register/C3689  ( .a(\prgm_register/en_not ), .b(a[202]), .out(
        \prgm_register/n406 ) );
  nand2 \prgm_register/C3690  ( .a(\prgm_register/n405 ), .b(
        \prgm_register/n406 ), .out(\prgm_register/or_signal [202]) );
  nand2 \prgm_register/C3691  ( .a(enable), .b(a[202]), .out(
        \prgm_register/n407 ) );
  nand2 \prgm_register/C3692  ( .a(\prgm_register/en_not ), .b(a[203]), .out(
        \prgm_register/n408 ) );
  nand2 \prgm_register/C3693  ( .a(\prgm_register/n407 ), .b(
        \prgm_register/n408 ), .out(\prgm_register/or_signal [203]) );
  nand2 \prgm_register/C3694  ( .a(enable), .b(a[203]), .out(
        \prgm_register/n409 ) );
  nand2 \prgm_register/C3695  ( .a(\prgm_register/en_not ), .b(a[204]), .out(
        \prgm_register/n410 ) );
  nand2 \prgm_register/C3696  ( .a(\prgm_register/n409 ), .b(
        \prgm_register/n410 ), .out(\prgm_register/or_signal [204]) );
  nand2 \prgm_register/C3697  ( .a(enable), .b(a[204]), .out(
        \prgm_register/n411 ) );
  nand2 \prgm_register/C3698  ( .a(\prgm_register/en_not ), .b(a[205]), .out(
        \prgm_register/n412 ) );
  nand2 \prgm_register/C3699  ( .a(\prgm_register/n411 ), .b(
        \prgm_register/n412 ), .out(\prgm_register/or_signal [205]) );
  nand2 \prgm_register/C3700  ( .a(enable), .b(a[205]), .out(
        \prgm_register/n413 ) );
  nand2 \prgm_register/C3701  ( .a(\prgm_register/en_not ), .b(a[206]), .out(
        \prgm_register/n414 ) );
  nand2 \prgm_register/C3702  ( .a(\prgm_register/n413 ), .b(
        \prgm_register/n414 ), .out(\prgm_register/or_signal [206]) );
  nand2 \prgm_register/C3703  ( .a(enable), .b(a[206]), .out(
        \prgm_register/n415 ) );
  nand2 \prgm_register/C3704  ( .a(\prgm_register/en_not ), .b(a[207]), .out(
        \prgm_register/n416 ) );
  nand2 \prgm_register/C3705  ( .a(\prgm_register/n415 ), .b(
        \prgm_register/n416 ), .out(\prgm_register/or_signal [207]) );
  nand2 \prgm_register/C3706  ( .a(enable), .b(a[207]), .out(
        \prgm_register/n417 ) );
  nand2 \prgm_register/C3707  ( .a(\prgm_register/en_not ), .b(a[208]), .out(
        \prgm_register/n418 ) );
  nand2 \prgm_register/C3708  ( .a(\prgm_register/n417 ), .b(
        \prgm_register/n418 ), .out(\prgm_register/or_signal [208]) );
  nand2 \prgm_register/C3709  ( .a(enable), .b(a[208]), .out(
        \prgm_register/n419 ) );
  nand2 \prgm_register/C3710  ( .a(\prgm_register/en_not ), .b(a[209]), .out(
        \prgm_register/n420 ) );
  nand2 \prgm_register/C3711  ( .a(\prgm_register/n419 ), .b(
        \prgm_register/n420 ), .out(\prgm_register/or_signal [209]) );
  nand2 \prgm_register/C3712  ( .a(enable), .b(a[209]), .out(
        \prgm_register/n421 ) );
  nand2 \prgm_register/C3713  ( .a(\prgm_register/en_not ), .b(a[210]), .out(
        \prgm_register/n422 ) );
  nand2 \prgm_register/C3714  ( .a(\prgm_register/n421 ), .b(
        \prgm_register/n422 ), .out(\prgm_register/or_signal [210]) );
  nand2 \prgm_register/C3715  ( .a(enable), .b(a[210]), .out(
        \prgm_register/n423 ) );
  nand2 \prgm_register/C3716  ( .a(\prgm_register/en_not ), .b(a[211]), .out(
        \prgm_register/n424 ) );
  nand2 \prgm_register/C3717  ( .a(\prgm_register/n423 ), .b(
        \prgm_register/n424 ), .out(\prgm_register/or_signal [211]) );
  nand2 \prgm_register/C3718  ( .a(enable), .b(a[211]), .out(
        \prgm_register/n425 ) );
  nand2 \prgm_register/C3719  ( .a(\prgm_register/en_not ), .b(a[212]), .out(
        \prgm_register/n426 ) );
  nand2 \prgm_register/C3720  ( .a(\prgm_register/n425 ), .b(
        \prgm_register/n426 ), .out(\prgm_register/or_signal [212]) );
  nand2 \prgm_register/C3721  ( .a(enable), .b(a[212]), .out(
        \prgm_register/n427 ) );
  nand2 \prgm_register/C3722  ( .a(\prgm_register/en_not ), .b(a[213]), .out(
        \prgm_register/n428 ) );
  nand2 \prgm_register/C3723  ( .a(\prgm_register/n427 ), .b(
        \prgm_register/n428 ), .out(\prgm_register/or_signal [213]) );
  nand2 \prgm_register/C3724  ( .a(enable), .b(a[213]), .out(
        \prgm_register/n429 ) );
  nand2 \prgm_register/C3725  ( .a(\prgm_register/en_not ), .b(a[214]), .out(
        \prgm_register/n430 ) );
  nand2 \prgm_register/C3726  ( .a(\prgm_register/n429 ), .b(
        \prgm_register/n430 ), .out(\prgm_register/or_signal [214]) );
  nand2 \prgm_register/C3727  ( .a(enable), .b(a[214]), .out(
        \prgm_register/n431 ) );
  nand2 \prgm_register/C3728  ( .a(\prgm_register/en_not ), .b(a[215]), .out(
        \prgm_register/n432 ) );
  nand2 \prgm_register/C3729  ( .a(\prgm_register/n431 ), .b(
        \prgm_register/n432 ), .out(\prgm_register/or_signal [215]) );
  nand2 \prgm_register/C3730  ( .a(enable), .b(a[215]), .out(
        \prgm_register/n433 ) );
  nand2 \prgm_register/C3731  ( .a(\prgm_register/en_not ), .b(a[216]), .out(
        \prgm_register/n434 ) );
  nand2 \prgm_register/C3732  ( .a(\prgm_register/n433 ), .b(
        \prgm_register/n434 ), .out(\prgm_register/or_signal [216]) );
  nand2 \prgm_register/C3733  ( .a(enable), .b(a[216]), .out(
        \prgm_register/n435 ) );
  nand2 \prgm_register/C3734  ( .a(\prgm_register/en_not ), .b(a[217]), .out(
        \prgm_register/n436 ) );
  nand2 \prgm_register/C3735  ( .a(\prgm_register/n435 ), .b(
        \prgm_register/n436 ), .out(\prgm_register/or_signal [217]) );
  nand2 \prgm_register/C3736  ( .a(enable), .b(a[217]), .out(
        \prgm_register/n437 ) );
  nand2 \prgm_register/C3737  ( .a(\prgm_register/en_not ), .b(a[218]), .out(
        \prgm_register/n438 ) );
  nand2 \prgm_register/C3738  ( .a(\prgm_register/n437 ), .b(
        \prgm_register/n438 ), .out(\prgm_register/or_signal [218]) );
  nand2 \prgm_register/C3739  ( .a(enable), .b(a[218]), .out(
        \prgm_register/n439 ) );
  nand2 \prgm_register/C3740  ( .a(\prgm_register/en_not ), .b(a[219]), .out(
        \prgm_register/n440 ) );
  nand2 \prgm_register/C3741  ( .a(\prgm_register/n439 ), .b(
        \prgm_register/n440 ), .out(\prgm_register/or_signal [219]) );
  nand2 \prgm_register/C3742  ( .a(enable), .b(a[219]), .out(
        \prgm_register/n441 ) );
  nand2 \prgm_register/C3743  ( .a(\prgm_register/en_not ), .b(a[220]), .out(
        \prgm_register/n442 ) );
  nand2 \prgm_register/C3744  ( .a(\prgm_register/n441 ), .b(
        \prgm_register/n442 ), .out(\prgm_register/or_signal [220]) );
  nand2 \prgm_register/C3745  ( .a(enable), .b(a[220]), .out(
        \prgm_register/n443 ) );
  nand2 \prgm_register/C3746  ( .a(\prgm_register/en_not ), .b(a[221]), .out(
        \prgm_register/n444 ) );
  nand2 \prgm_register/C3747  ( .a(\prgm_register/n443 ), .b(
        \prgm_register/n444 ), .out(\prgm_register/or_signal [221]) );
  nand2 \prgm_register/C3748  ( .a(enable), .b(a[221]), .out(
        \prgm_register/n445 ) );
  nand2 \prgm_register/C3749  ( .a(\prgm_register/en_not ), .b(a[222]), .out(
        \prgm_register/n446 ) );
  nand2 \prgm_register/C3750  ( .a(\prgm_register/n445 ), .b(
        \prgm_register/n446 ), .out(\prgm_register/or_signal [222]) );
  nand2 \prgm_register/C3751  ( .a(enable), .b(a[222]), .out(
        \prgm_register/n447 ) );
  nand2 \prgm_register/C3752  ( .a(\prgm_register/en_not ), .b(a[223]), .out(
        \prgm_register/n448 ) );
  nand2 \prgm_register/C3753  ( .a(\prgm_register/n447 ), .b(
        \prgm_register/n448 ), .out(\prgm_register/or_signal [223]) );
  nand2 \prgm_register/C3754  ( .a(enable), .b(a[223]), .out(
        \prgm_register/n449 ) );
  nand2 \prgm_register/C3755  ( .a(\prgm_register/en_not ), .b(a[224]), .out(
        \prgm_register/n450 ) );
  nand2 \prgm_register/C3756  ( .a(\prgm_register/n449 ), .b(
        \prgm_register/n450 ), .out(\prgm_register/or_signal [224]) );
  nand2 \prgm_register/C3757  ( .a(enable), .b(a[224]), .out(
        \prgm_register/n451 ) );
  nand2 \prgm_register/C3758  ( .a(\prgm_register/en_not ), .b(a[225]), .out(
        \prgm_register/n452 ) );
  nand2 \prgm_register/C3759  ( .a(\prgm_register/n451 ), .b(
        \prgm_register/n452 ), .out(\prgm_register/or_signal [225]) );
  nand2 \prgm_register/C3760  ( .a(enable), .b(a[225]), .out(
        \prgm_register/n453 ) );
  nand2 \prgm_register/C3761  ( .a(\prgm_register/en_not ), .b(a[226]), .out(
        \prgm_register/n454 ) );
  nand2 \prgm_register/C3762  ( .a(\prgm_register/n453 ), .b(
        \prgm_register/n454 ), .out(\prgm_register/or_signal [226]) );
  nand2 \prgm_register/C3763  ( .a(enable), .b(a[226]), .out(
        \prgm_register/n455 ) );
  nand2 \prgm_register/C3764  ( .a(\prgm_register/en_not ), .b(a[227]), .out(
        \prgm_register/n456 ) );
  nand2 \prgm_register/C3765  ( .a(\prgm_register/n455 ), .b(
        \prgm_register/n456 ), .out(\prgm_register/or_signal [227]) );
  nand2 \prgm_register/C3766  ( .a(enable), .b(a[227]), .out(
        \prgm_register/n457 ) );
  nand2 \prgm_register/C3767  ( .a(\prgm_register/en_not ), .b(a[228]), .out(
        \prgm_register/n458 ) );
  nand2 \prgm_register/C3768  ( .a(\prgm_register/n457 ), .b(
        \prgm_register/n458 ), .out(\prgm_register/or_signal [228]) );
  nand2 \prgm_register/C3769  ( .a(enable), .b(a[228]), .out(
        \prgm_register/n459 ) );
  nand2 \prgm_register/C3770  ( .a(\prgm_register/en_not ), .b(a[229]), .out(
        \prgm_register/n460 ) );
  nand2 \prgm_register/C3771  ( .a(\prgm_register/n459 ), .b(
        \prgm_register/n460 ), .out(\prgm_register/or_signal [229]) );
  nand2 \prgm_register/C3772  ( .a(enable), .b(a[229]), .out(
        \prgm_register/n461 ) );
  nand2 \prgm_register/C3773  ( .a(\prgm_register/en_not ), .b(a[230]), .out(
        \prgm_register/n462 ) );
  nand2 \prgm_register/C3774  ( .a(\prgm_register/n461 ), .b(
        \prgm_register/n462 ), .out(\prgm_register/or_signal [230]) );
  nand2 \prgm_register/C3775  ( .a(enable), .b(a[230]), .out(
        \prgm_register/n463 ) );
  nand2 \prgm_register/C3776  ( .a(\prgm_register/en_not ), .b(a[231]), .out(
        \prgm_register/n464 ) );
  nand2 \prgm_register/C3777  ( .a(\prgm_register/n463 ), .b(
        \prgm_register/n464 ), .out(\prgm_register/or_signal [231]) );
  nand2 \prgm_register/C3778  ( .a(enable), .b(a[231]), .out(
        \prgm_register/n465 ) );
  nand2 \prgm_register/C3779  ( .a(\prgm_register/en_not ), .b(a[232]), .out(
        \prgm_register/n466 ) );
  nand2 \prgm_register/C3780  ( .a(\prgm_register/n465 ), .b(
        \prgm_register/n466 ), .out(\prgm_register/or_signal [232]) );
  nand2 \prgm_register/C3781  ( .a(enable), .b(a[232]), .out(
        \prgm_register/n467 ) );
  nand2 \prgm_register/C3782  ( .a(\prgm_register/en_not ), .b(a[233]), .out(
        \prgm_register/n468 ) );
  nand2 \prgm_register/C3783  ( .a(\prgm_register/n467 ), .b(
        \prgm_register/n468 ), .out(\prgm_register/or_signal [233]) );
  nand2 \prgm_register/C3784  ( .a(enable), .b(a[233]), .out(
        \prgm_register/n469 ) );
  nand2 \prgm_register/C3785  ( .a(\prgm_register/en_not ), .b(a[234]), .out(
        \prgm_register/n470 ) );
  nand2 \prgm_register/C3786  ( .a(\prgm_register/n469 ), .b(
        \prgm_register/n470 ), .out(\prgm_register/or_signal [234]) );
  nand2 \prgm_register/C3787  ( .a(enable), .b(a[234]), .out(
        \prgm_register/n471 ) );
  nand2 \prgm_register/C3788  ( .a(\prgm_register/en_not ), .b(a[235]), .out(
        \prgm_register/n472 ) );
  nand2 \prgm_register/C3789  ( .a(\prgm_register/n471 ), .b(
        \prgm_register/n472 ), .out(\prgm_register/or_signal [235]) );
  nand2 \prgm_register/C3790  ( .a(enable), .b(a[235]), .out(
        \prgm_register/n473 ) );
  nand2 \prgm_register/C3791  ( .a(\prgm_register/en_not ), .b(a[236]), .out(
        \prgm_register/n474 ) );
  nand2 \prgm_register/C3792  ( .a(\prgm_register/n473 ), .b(
        \prgm_register/n474 ), .out(\prgm_register/or_signal [236]) );
  nand2 \prgm_register/C3793  ( .a(enable), .b(a[236]), .out(
        \prgm_register/n475 ) );
  nand2 \prgm_register/C3794  ( .a(\prgm_register/en_not ), .b(a[237]), .out(
        \prgm_register/n476 ) );
  nand2 \prgm_register/C3795  ( .a(\prgm_register/n475 ), .b(
        \prgm_register/n476 ), .out(\prgm_register/or_signal [237]) );
  nand2 \prgm_register/C3796  ( .a(enable), .b(a[237]), .out(
        \prgm_register/n477 ) );
  nand2 \prgm_register/C3797  ( .a(\prgm_register/en_not ), .b(a[238]), .out(
        \prgm_register/n478 ) );
  nand2 \prgm_register/C3798  ( .a(\prgm_register/n477 ), .b(
        \prgm_register/n478 ), .out(\prgm_register/or_signal [238]) );
  nand2 \prgm_register/C3799  ( .a(enable), .b(a[238]), .out(
        \prgm_register/n479 ) );
  nand2 \prgm_register/C3800  ( .a(\prgm_register/en_not ), .b(a[239]), .out(
        \prgm_register/n480 ) );
  nand2 \prgm_register/C3801  ( .a(\prgm_register/n479 ), .b(
        \prgm_register/n480 ), .out(\prgm_register/or_signal [239]) );
  nand2 \prgm_register/C3802  ( .a(enable), .b(a[239]), .out(
        \prgm_register/n481 ) );
  nand2 \prgm_register/C3803  ( .a(\prgm_register/en_not ), .b(a[240]), .out(
        \prgm_register/n482 ) );
  nand2 \prgm_register/C3804  ( .a(\prgm_register/n481 ), .b(
        \prgm_register/n482 ), .out(\prgm_register/or_signal [240]) );
  nand2 \prgm_register/C3805  ( .a(enable), .b(a[240]), .out(
        \prgm_register/n483 ) );
  nand2 \prgm_register/C3806  ( .a(\prgm_register/en_not ), .b(a[241]), .out(
        \prgm_register/n484 ) );
  nand2 \prgm_register/C3807  ( .a(\prgm_register/n483 ), .b(
        \prgm_register/n484 ), .out(\prgm_register/or_signal [241]) );
  nand2 \prgm_register/C3808  ( .a(enable), .b(a[241]), .out(
        \prgm_register/n485 ) );
  nand2 \prgm_register/C3809  ( .a(\prgm_register/en_not ), .b(a[242]), .out(
        \prgm_register/n486 ) );
  nand2 \prgm_register/C3810  ( .a(\prgm_register/n485 ), .b(
        \prgm_register/n486 ), .out(\prgm_register/or_signal [242]) );
  nand2 \prgm_register/C3811  ( .a(enable), .b(a[242]), .out(
        \prgm_register/n487 ) );
  nand2 \prgm_register/C3812  ( .a(\prgm_register/en_not ), .b(a[243]), .out(
        \prgm_register/n488 ) );
  nand2 \prgm_register/C3813  ( .a(\prgm_register/n487 ), .b(
        \prgm_register/n488 ), .out(\prgm_register/or_signal [243]) );
  nand2 \prgm_register/C3814  ( .a(enable), .b(a[243]), .out(
        \prgm_register/n489 ) );
  nand2 \prgm_register/C3815  ( .a(\prgm_register/en_not ), .b(a[244]), .out(
        \prgm_register/n490 ) );
  nand2 \prgm_register/C3816  ( .a(\prgm_register/n489 ), .b(
        \prgm_register/n490 ), .out(\prgm_register/or_signal [244]) );
  nand2 \prgm_register/C3817  ( .a(enable), .b(a[244]), .out(
        \prgm_register/n491 ) );
  nand2 \prgm_register/C3818  ( .a(\prgm_register/en_not ), .b(a[245]), .out(
        \prgm_register/n492 ) );
  nand2 \prgm_register/C3819  ( .a(\prgm_register/n491 ), .b(
        \prgm_register/n492 ), .out(\prgm_register/or_signal [245]) );
  nand2 \prgm_register/C3820  ( .a(enable), .b(a[245]), .out(
        \prgm_register/n493 ) );
  nand2 \prgm_register/C3821  ( .a(\prgm_register/en_not ), .b(a[246]), .out(
        \prgm_register/n494 ) );
  nand2 \prgm_register/C3822  ( .a(\prgm_register/n493 ), .b(
        \prgm_register/n494 ), .out(\prgm_register/or_signal [246]) );
  nand2 \prgm_register/C3823  ( .a(enable), .b(a[246]), .out(
        \prgm_register/n495 ) );
  nand2 \prgm_register/C3824  ( .a(\prgm_register/en_not ), .b(a[247]), .out(
        \prgm_register/n496 ) );
  nand2 \prgm_register/C3825  ( .a(\prgm_register/n495 ), .b(
        \prgm_register/n496 ), .out(\prgm_register/or_signal [247]) );
  nand2 \prgm_register/C3826  ( .a(enable), .b(a[247]), .out(
        \prgm_register/n497 ) );
  nand2 \prgm_register/C3827  ( .a(\prgm_register/en_not ), .b(a[248]), .out(
        \prgm_register/n498 ) );
  nand2 \prgm_register/C3828  ( .a(\prgm_register/n497 ), .b(
        \prgm_register/n498 ), .out(\prgm_register/or_signal [248]) );
  nand2 \prgm_register/C3829  ( .a(enable), .b(a[248]), .out(
        \prgm_register/n499 ) );
  nand2 \prgm_register/C3830  ( .a(\prgm_register/en_not ), .b(a[249]), .out(
        \prgm_register/n500 ) );
  nand2 \prgm_register/C3831  ( .a(\prgm_register/n499 ), .b(
        \prgm_register/n500 ), .out(\prgm_register/or_signal [249]) );
  nand2 \prgm_register/C3832  ( .a(enable), .b(a[249]), .out(
        \prgm_register/n501 ) );
  nand2 \prgm_register/C3833  ( .a(\prgm_register/en_not ), .b(a[250]), .out(
        \prgm_register/n502 ) );
  nand2 \prgm_register/C3834  ( .a(\prgm_register/n501 ), .b(
        \prgm_register/n502 ), .out(\prgm_register/or_signal [250]) );
  nand2 \prgm_register/C3835  ( .a(enable), .b(a[250]), .out(
        \prgm_register/n503 ) );
  nand2 \prgm_register/C3836  ( .a(\prgm_register/en_not ), .b(a[251]), .out(
        \prgm_register/n504 ) );
  nand2 \prgm_register/C3837  ( .a(\prgm_register/n503 ), .b(
        \prgm_register/n504 ), .out(\prgm_register/or_signal [251]) );
  nand2 \prgm_register/C3838  ( .a(enable), .b(a[251]), .out(
        \prgm_register/n505 ) );
  nand2 \prgm_register/C3839  ( .a(\prgm_register/en_not ), .b(a[252]), .out(
        \prgm_register/n506 ) );
  nand2 \prgm_register/C3840  ( .a(\prgm_register/n505 ), .b(
        \prgm_register/n506 ), .out(\prgm_register/or_signal [252]) );
  nand2 \prgm_register/C3841  ( .a(enable), .b(a[252]), .out(
        \prgm_register/n507 ) );
  nand2 \prgm_register/C3842  ( .a(\prgm_register/en_not ), .b(a[253]), .out(
        \prgm_register/n508 ) );
  nand2 \prgm_register/C3843  ( .a(\prgm_register/n507 ), .b(
        \prgm_register/n508 ), .out(\prgm_register/or_signal [253]) );
  nand2 \prgm_register/C3844  ( .a(enable), .b(a[253]), .out(
        \prgm_register/n509 ) );
  nand2 \prgm_register/C3845  ( .a(\prgm_register/en_not ), .b(a[254]), .out(
        \prgm_register/n510 ) );
  nand2 \prgm_register/C3846  ( .a(\prgm_register/n509 ), .b(
        \prgm_register/n510 ), .out(\prgm_register/or_signal [254]) );
  nand2 \prgm_register/C3847  ( .a(enable), .b(a[254]), .out(
        \prgm_register/n511 ) );
  nand2 \prgm_register/C3848  ( .a(\prgm_register/en_not ), .b(a[255]), .out(
        \prgm_register/n512 ) );
  nand2 \prgm_register/C3849  ( .a(\prgm_register/n511 ), .b(
        \prgm_register/n512 ), .out(\prgm_register/or_signal [255]) );
  nand2 \prgm_register/C3850  ( .a(enable), .b(a[255]), .out(
        \prgm_register/n513 ) );
  nand2 \prgm_register/C3851  ( .a(\prgm_register/en_not ), .b(a[256]), .out(
        \prgm_register/n514 ) );
  nand2 \prgm_register/C3852  ( .a(\prgm_register/n513 ), .b(
        \prgm_register/n514 ), .out(\prgm_register/or_signal [256]) );
  nand2 \prgm_register/C3853  ( .a(enable), .b(a[256]), .out(
        \prgm_register/n515 ) );
  nand2 \prgm_register/C3854  ( .a(\prgm_register/en_not ), .b(a[257]), .out(
        \prgm_register/n516 ) );
  nand2 \prgm_register/C3855  ( .a(\prgm_register/n515 ), .b(
        \prgm_register/n516 ), .out(\prgm_register/or_signal [257]) );
  nand2 \prgm_register/C3856  ( .a(enable), .b(a[257]), .out(
        \prgm_register/n517 ) );
  nand2 \prgm_register/C3857  ( .a(\prgm_register/en_not ), .b(a[258]), .out(
        \prgm_register/n518 ) );
  nand2 \prgm_register/C3858  ( .a(\prgm_register/n517 ), .b(
        \prgm_register/n518 ), .out(\prgm_register/or_signal [258]) );
  nand2 \prgm_register/C3859  ( .a(enable), .b(a[258]), .out(
        \prgm_register/n519 ) );
  nand2 \prgm_register/C3860  ( .a(\prgm_register/en_not ), .b(a[259]), .out(
        \prgm_register/n520 ) );
  nand2 \prgm_register/C3861  ( .a(\prgm_register/n519 ), .b(
        \prgm_register/n520 ), .out(\prgm_register/or_signal [259]) );
  nand2 \prgm_register/C3862  ( .a(enable), .b(a[259]), .out(
        \prgm_register/n521 ) );
  nand2 \prgm_register/C3863  ( .a(\prgm_register/en_not ), .b(a[260]), .out(
        \prgm_register/n522 ) );
  nand2 \prgm_register/C3864  ( .a(\prgm_register/n521 ), .b(
        \prgm_register/n522 ), .out(\prgm_register/or_signal [260]) );
  nand2 \prgm_register/C3865  ( .a(enable), .b(a[260]), .out(
        \prgm_register/n523 ) );
  nand2 \prgm_register/C3866  ( .a(\prgm_register/en_not ), .b(a[261]), .out(
        \prgm_register/n524 ) );
  nand2 \prgm_register/C3867  ( .a(\prgm_register/n523 ), .b(
        \prgm_register/n524 ), .out(\prgm_register/or_signal [261]) );
  nand2 \prgm_register/C3868  ( .a(enable), .b(a[261]), .out(
        \prgm_register/n525 ) );
  nand2 \prgm_register/C3869  ( .a(\prgm_register/en_not ), .b(a[262]), .out(
        \prgm_register/n526 ) );
  nand2 \prgm_register/C3870  ( .a(\prgm_register/n525 ), .b(
        \prgm_register/n526 ), .out(\prgm_register/or_signal [262]) );
  nand2 \prgm_register/C3871  ( .a(enable), .b(a[262]), .out(
        \prgm_register/n527 ) );
  nand2 \prgm_register/C3872  ( .a(\prgm_register/en_not ), .b(a[263]), .out(
        \prgm_register/n528 ) );
  nand2 \prgm_register/C3873  ( .a(\prgm_register/n527 ), .b(
        \prgm_register/n528 ), .out(\prgm_register/or_signal [263]) );
  nand2 \prgm_register/C3874  ( .a(enable), .b(a[263]), .out(
        \prgm_register/n529 ) );
  nand2 \prgm_register/C3875  ( .a(\prgm_register/en_not ), .b(a[264]), .out(
        \prgm_register/n530 ) );
  nand2 \prgm_register/C3876  ( .a(\prgm_register/n529 ), .b(
        \prgm_register/n530 ), .out(\prgm_register/or_signal [264]) );
  nand2 \prgm_register/C3877  ( .a(enable), .b(a[264]), .out(
        \prgm_register/n531 ) );
  nand2 \prgm_register/C3878  ( .a(\prgm_register/en_not ), .b(a[265]), .out(
        \prgm_register/n532 ) );
  nand2 \prgm_register/C3879  ( .a(\prgm_register/n531 ), .b(
        \prgm_register/n532 ), .out(\prgm_register/or_signal [265]) );
  nand2 \prgm_register/C3880  ( .a(enable), .b(a[265]), .out(
        \prgm_register/n533 ) );
  nand2 \prgm_register/C3881  ( .a(\prgm_register/en_not ), .b(a[266]), .out(
        \prgm_register/n534 ) );
  nand2 \prgm_register/C3882  ( .a(\prgm_register/n533 ), .b(
        \prgm_register/n534 ), .out(\prgm_register/or_signal [266]) );
  nand2 \prgm_register/C3883  ( .a(enable), .b(a[266]), .out(
        \prgm_register/n535 ) );
  nand2 \prgm_register/C3884  ( .a(\prgm_register/en_not ), .b(a[267]), .out(
        \prgm_register/n536 ) );
  nand2 \prgm_register/C3885  ( .a(\prgm_register/n535 ), .b(
        \prgm_register/n536 ), .out(\prgm_register/or_signal [267]) );
  nand2 \prgm_register/C3886  ( .a(enable), .b(a[267]), .out(
        \prgm_register/n537 ) );
  nand2 \prgm_register/C3887  ( .a(\prgm_register/en_not ), .b(a[268]), .out(
        \prgm_register/n538 ) );
  nand2 \prgm_register/C3888  ( .a(\prgm_register/n537 ), .b(
        \prgm_register/n538 ), .out(\prgm_register/or_signal [268]) );
  nand2 \prgm_register/C3889  ( .a(enable), .b(a[268]), .out(
        \prgm_register/n539 ) );
  nand2 \prgm_register/C3890  ( .a(\prgm_register/en_not ), .b(a[269]), .out(
        \prgm_register/n540 ) );
  nand2 \prgm_register/C3891  ( .a(\prgm_register/n539 ), .b(
        \prgm_register/n540 ), .out(\prgm_register/or_signal [269]) );
  nand2 \prgm_register/C3892  ( .a(enable), .b(a[269]), .out(
        \prgm_register/n541 ) );
  nand2 \prgm_register/C3893  ( .a(\prgm_register/en_not ), .b(a[270]), .out(
        \prgm_register/n542 ) );
  nand2 \prgm_register/C3894  ( .a(\prgm_register/n541 ), .b(
        \prgm_register/n542 ), .out(\prgm_register/or_signal [270]) );
  nand2 \prgm_register/C3895  ( .a(enable), .b(a[270]), .out(
        \prgm_register/n543 ) );
  nand2 \prgm_register/C3896  ( .a(\prgm_register/en_not ), .b(a[271]), .out(
        \prgm_register/n544 ) );
  nand2 \prgm_register/C3897  ( .a(\prgm_register/n543 ), .b(
        \prgm_register/n544 ), .out(\prgm_register/or_signal [271]) );
  nand2 \prgm_register/C3898  ( .a(enable), .b(a[271]), .out(
        \prgm_register/n545 ) );
  nand2 \prgm_register/C3899  ( .a(\prgm_register/en_not ), .b(a[272]), .out(
        \prgm_register/n546 ) );
  nand2 \prgm_register/C3900  ( .a(\prgm_register/n545 ), .b(
        \prgm_register/n546 ), .out(\prgm_register/or_signal [272]) );
  nand2 \prgm_register/C3901  ( .a(enable), .b(a[272]), .out(
        \prgm_register/n547 ) );
  nand2 \prgm_register/C3902  ( .a(\prgm_register/en_not ), .b(a[273]), .out(
        \prgm_register/n548 ) );
  nand2 \prgm_register/C3903  ( .a(\prgm_register/n547 ), .b(
        \prgm_register/n548 ), .out(\prgm_register/or_signal [273]) );
  nand2 \prgm_register/C3904  ( .a(enable), .b(a[273]), .out(
        \prgm_register/n549 ) );
  nand2 \prgm_register/C3905  ( .a(\prgm_register/en_not ), .b(a[274]), .out(
        \prgm_register/n550 ) );
  nand2 \prgm_register/C3906  ( .a(\prgm_register/n549 ), .b(
        \prgm_register/n550 ), .out(\prgm_register/or_signal [274]) );
  nand2 \prgm_register/C3907  ( .a(enable), .b(a[274]), .out(
        \prgm_register/n551 ) );
  nand2 \prgm_register/C3908  ( .a(\prgm_register/en_not ), .b(a[275]), .out(
        \prgm_register/n552 ) );
  nand2 \prgm_register/C3909  ( .a(\prgm_register/n551 ), .b(
        \prgm_register/n552 ), .out(\prgm_register/or_signal [275]) );
  nand2 \prgm_register/C3910  ( .a(enable), .b(a[275]), .out(
        \prgm_register/n553 ) );
  nand2 \prgm_register/C3911  ( .a(\prgm_register/en_not ), .b(a[276]), .out(
        \prgm_register/n554 ) );
  nand2 \prgm_register/C3912  ( .a(\prgm_register/n553 ), .b(
        \prgm_register/n554 ), .out(\prgm_register/or_signal [276]) );
  nand2 \prgm_register/C3913  ( .a(enable), .b(a[276]), .out(
        \prgm_register/n555 ) );
  nand2 \prgm_register/C3914  ( .a(\prgm_register/en_not ), .b(a[277]), .out(
        \prgm_register/n556 ) );
  nand2 \prgm_register/C3915  ( .a(\prgm_register/n555 ), .b(
        \prgm_register/n556 ), .out(\prgm_register/or_signal [277]) );
  nand2 \prgm_register/C3916  ( .a(enable), .b(a[277]), .out(
        \prgm_register/n557 ) );
  nand2 \prgm_register/C3917  ( .a(\prgm_register/en_not ), .b(a[278]), .out(
        \prgm_register/n558 ) );
  nand2 \prgm_register/C3918  ( .a(\prgm_register/n557 ), .b(
        \prgm_register/n558 ), .out(\prgm_register/or_signal [278]) );
  nand2 \prgm_register/C3919  ( .a(enable), .b(a[278]), .out(
        \prgm_register/n559 ) );
  nand2 \prgm_register/C3920  ( .a(\prgm_register/en_not ), .b(a[279]), .out(
        \prgm_register/n560 ) );
  nand2 \prgm_register/C3921  ( .a(\prgm_register/n559 ), .b(
        \prgm_register/n560 ), .out(\prgm_register/or_signal [279]) );
  nand2 \prgm_register/C3922  ( .a(enable), .b(a[279]), .out(
        \prgm_register/n561 ) );
  nand2 \prgm_register/C3923  ( .a(\prgm_register/en_not ), .b(a[280]), .out(
        \prgm_register/n562 ) );
  nand2 \prgm_register/C3924  ( .a(\prgm_register/n561 ), .b(
        \prgm_register/n562 ), .out(\prgm_register/or_signal [280]) );
  nand2 \prgm_register/C3925  ( .a(enable), .b(a[280]), .out(
        \prgm_register/n563 ) );
  nand2 \prgm_register/C3926  ( .a(\prgm_register/en_not ), .b(a[281]), .out(
        \prgm_register/n564 ) );
  nand2 \prgm_register/C3927  ( .a(\prgm_register/n563 ), .b(
        \prgm_register/n564 ), .out(\prgm_register/or_signal [281]) );
  nand2 \prgm_register/C3928  ( .a(enable), .b(a[281]), .out(
        \prgm_register/n565 ) );
  nand2 \prgm_register/C3929  ( .a(\prgm_register/en_not ), .b(a[282]), .out(
        \prgm_register/n566 ) );
  nand2 \prgm_register/C3930  ( .a(\prgm_register/n565 ), .b(
        \prgm_register/n566 ), .out(\prgm_register/or_signal [282]) );
  nand2 \prgm_register/C3931  ( .a(enable), .b(a[282]), .out(
        \prgm_register/n567 ) );
  nand2 \prgm_register/C3932  ( .a(\prgm_register/en_not ), .b(a[283]), .out(
        \prgm_register/n568 ) );
  nand2 \prgm_register/C3933  ( .a(\prgm_register/n567 ), .b(
        \prgm_register/n568 ), .out(\prgm_register/or_signal [283]) );
  nand2 \prgm_register/C3934  ( .a(enable), .b(a[283]), .out(
        \prgm_register/n569 ) );
  nand2 \prgm_register/C3935  ( .a(\prgm_register/en_not ), .b(a[284]), .out(
        \prgm_register/n570 ) );
  nand2 \prgm_register/C3936  ( .a(\prgm_register/n569 ), .b(
        \prgm_register/n570 ), .out(\prgm_register/or_signal [284]) );
  nand2 \prgm_register/C3937  ( .a(enable), .b(a[284]), .out(
        \prgm_register/n571 ) );
  nand2 \prgm_register/C3938  ( .a(\prgm_register/en_not ), .b(a[285]), .out(
        \prgm_register/n572 ) );
  nand2 \prgm_register/C3939  ( .a(\prgm_register/n571 ), .b(
        \prgm_register/n572 ), .out(\prgm_register/or_signal [285]) );
  nand2 \prgm_register/C3940  ( .a(enable), .b(a[285]), .out(
        \prgm_register/n573 ) );
  nand2 \prgm_register/C3941  ( .a(\prgm_register/en_not ), .b(a[286]), .out(
        \prgm_register/n574 ) );
  nand2 \prgm_register/C3942  ( .a(\prgm_register/n573 ), .b(
        \prgm_register/n574 ), .out(\prgm_register/or_signal [286]) );
  nand2 \prgm_register/C3943  ( .a(enable), .b(a[286]), .out(
        \prgm_register/n575 ) );
  nand2 \prgm_register/C3944  ( .a(\prgm_register/en_not ), .b(a[287]), .out(
        \prgm_register/n576 ) );
  nand2 \prgm_register/C3945  ( .a(\prgm_register/n575 ), .b(
        \prgm_register/n576 ), .out(\prgm_register/or_signal [287]) );
  nand2 \prgm_register/C3946  ( .a(enable), .b(a[287]), .out(
        \prgm_register/n577 ) );
  nand2 \prgm_register/C3947  ( .a(\prgm_register/en_not ), .b(a[288]), .out(
        \prgm_register/n578 ) );
  nand2 \prgm_register/C3948  ( .a(\prgm_register/n577 ), .b(
        \prgm_register/n578 ), .out(\prgm_register/or_signal [288]) );
  nand2 \prgm_register/C3949  ( .a(enable), .b(a[288]), .out(
        \prgm_register/n579 ) );
  nand2 \prgm_register/C3950  ( .a(\prgm_register/en_not ), .b(a[289]), .out(
        \prgm_register/n580 ) );
  nand2 \prgm_register/C3951  ( .a(\prgm_register/n579 ), .b(
        \prgm_register/n580 ), .out(\prgm_register/or_signal [289]) );
  nand2 \prgm_register/C3952  ( .a(enable), .b(a[289]), .out(
        \prgm_register/n581 ) );
  nand2 \prgm_register/C3953  ( .a(\prgm_register/en_not ), .b(a[290]), .out(
        \prgm_register/n582 ) );
  nand2 \prgm_register/C3954  ( .a(\prgm_register/n581 ), .b(
        \prgm_register/n582 ), .out(\prgm_register/or_signal [290]) );
  nand2 \prgm_register/C3955  ( .a(enable), .b(a[290]), .out(
        \prgm_register/n583 ) );
  nand2 \prgm_register/C3956  ( .a(\prgm_register/en_not ), .b(a[291]), .out(
        \prgm_register/n584 ) );
  nand2 \prgm_register/C3957  ( .a(\prgm_register/n583 ), .b(
        \prgm_register/n584 ), .out(\prgm_register/or_signal [291]) );
  nand2 \prgm_register/C3958  ( .a(enable), .b(a[291]), .out(
        \prgm_register/n585 ) );
  nand2 \prgm_register/C3959  ( .a(\prgm_register/en_not ), .b(a[292]), .out(
        \prgm_register/n586 ) );
  nand2 \prgm_register/C3960  ( .a(\prgm_register/n585 ), .b(
        \prgm_register/n586 ), .out(\prgm_register/or_signal [292]) );
  nand2 \prgm_register/C3961  ( .a(enable), .b(a[292]), .out(
        \prgm_register/n587 ) );
  nand2 \prgm_register/C3962  ( .a(\prgm_register/en_not ), .b(a[293]), .out(
        \prgm_register/n588 ) );
  nand2 \prgm_register/C3963  ( .a(\prgm_register/n587 ), .b(
        \prgm_register/n588 ), .out(\prgm_register/or_signal [293]) );
  nand2 \prgm_register/C3964  ( .a(enable), .b(a[293]), .out(
        \prgm_register/n589 ) );
  nand2 \prgm_register/C3965  ( .a(\prgm_register/en_not ), .b(a[294]), .out(
        \prgm_register/n590 ) );
  nand2 \prgm_register/C3966  ( .a(\prgm_register/n589 ), .b(
        \prgm_register/n590 ), .out(\prgm_register/or_signal [294]) );
  nand2 \prgm_register/C3967  ( .a(enable), .b(a[294]), .out(
        \prgm_register/n591 ) );
  nand2 \prgm_register/C3968  ( .a(\prgm_register/en_not ), .b(a[295]), .out(
        \prgm_register/n592 ) );
  nand2 \prgm_register/C3969  ( .a(\prgm_register/n591 ), .b(
        \prgm_register/n592 ), .out(\prgm_register/or_signal [295]) );
  nand2 \prgm_register/C3970  ( .a(enable), .b(a[295]), .out(
        \prgm_register/n593 ) );
  nand2 \prgm_register/C3971  ( .a(\prgm_register/en_not ), .b(a[296]), .out(
        \prgm_register/n594 ) );
  nand2 \prgm_register/C3972  ( .a(\prgm_register/n593 ), .b(
        \prgm_register/n594 ), .out(\prgm_register/or_signal [296]) );
  nand2 \prgm_register/C3973  ( .a(enable), .b(a[296]), .out(
        \prgm_register/n595 ) );
  nand2 \prgm_register/C3974  ( .a(\prgm_register/en_not ), .b(a[297]), .out(
        \prgm_register/n596 ) );
  nand2 \prgm_register/C3975  ( .a(\prgm_register/n595 ), .b(
        \prgm_register/n596 ), .out(\prgm_register/or_signal [297]) );
  nand2 \prgm_register/C3976  ( .a(enable), .b(a[297]), .out(
        \prgm_register/n597 ) );
  nand2 \prgm_register/C3977  ( .a(\prgm_register/en_not ), .b(a[298]), .out(
        \prgm_register/n598 ) );
  nand2 \prgm_register/C3978  ( .a(\prgm_register/n597 ), .b(
        \prgm_register/n598 ), .out(\prgm_register/or_signal [298]) );
  nand2 \prgm_register/C3979  ( .a(enable), .b(a[298]), .out(
        \prgm_register/n599 ) );
  nand2 \prgm_register/C3980  ( .a(\prgm_register/en_not ), .b(a[299]), .out(
        \prgm_register/n600 ) );
  nand2 \prgm_register/C3981  ( .a(\prgm_register/n599 ), .b(
        \prgm_register/n600 ), .out(\prgm_register/or_signal [299]) );
  nand2 \prgm_register/C3982  ( .a(enable), .b(a[299]), .out(
        \prgm_register/n601 ) );
  nand2 \prgm_register/C3983  ( .a(\prgm_register/en_not ), .b(a[300]), .out(
        \prgm_register/n602 ) );
  nand2 \prgm_register/C3984  ( .a(\prgm_register/n601 ), .b(
        \prgm_register/n602 ), .out(\prgm_register/or_signal [300]) );
  nand2 \prgm_register/C3985  ( .a(enable), .b(a[300]), .out(
        \prgm_register/n603 ) );
  nand2 \prgm_register/C3986  ( .a(\prgm_register/en_not ), .b(a[301]), .out(
        \prgm_register/n604 ) );
  nand2 \prgm_register/C3987  ( .a(\prgm_register/n603 ), .b(
        \prgm_register/n604 ), .out(\prgm_register/or_signal [301]) );
  nand2 \prgm_register/C3988  ( .a(enable), .b(a[301]), .out(
        \prgm_register/n605 ) );
  nand2 \prgm_register/C3989  ( .a(\prgm_register/en_not ), .b(a[302]), .out(
        \prgm_register/n606 ) );
  nand2 \prgm_register/C3990  ( .a(\prgm_register/n605 ), .b(
        \prgm_register/n606 ), .out(\prgm_register/or_signal [302]) );
  nand2 \prgm_register/C3991  ( .a(enable), .b(a[302]), .out(
        \prgm_register/n607 ) );
  nand2 \prgm_register/C3992  ( .a(\prgm_register/en_not ), .b(a[303]), .out(
        \prgm_register/n608 ) );
  nand2 \prgm_register/C3993  ( .a(\prgm_register/n607 ), .b(
        \prgm_register/n608 ), .out(\prgm_register/or_signal [303]) );
  nand2 \prgm_register/C3994  ( .a(enable), .b(a[303]), .out(
        \prgm_register/n609 ) );
  nand2 \prgm_register/C3995  ( .a(\prgm_register/en_not ), .b(a[304]), .out(
        \prgm_register/n610 ) );
  nand2 \prgm_register/C3996  ( .a(\prgm_register/n609 ), .b(
        \prgm_register/n610 ), .out(\prgm_register/or_signal [304]) );
  nand2 \prgm_register/C3997  ( .a(enable), .b(a[304]), .out(
        \prgm_register/n611 ) );
  nand2 \prgm_register/C3998  ( .a(\prgm_register/en_not ), .b(a[305]), .out(
        \prgm_register/n612 ) );
  nand2 \prgm_register/C3999  ( .a(\prgm_register/n611 ), .b(
        \prgm_register/n612 ), .out(\prgm_register/or_signal [305]) );
  nand2 \prgm_register/C4000  ( .a(enable), .b(a[305]), .out(
        \prgm_register/n613 ) );
  nand2 \prgm_register/C4001  ( .a(\prgm_register/en_not ), .b(a[306]), .out(
        \prgm_register/n614 ) );
  nand2 \prgm_register/C4002  ( .a(\prgm_register/n613 ), .b(
        \prgm_register/n614 ), .out(\prgm_register/or_signal [306]) );
  nand2 \prgm_register/C4003  ( .a(enable), .b(a[306]), .out(
        \prgm_register/n615 ) );
  nand2 \prgm_register/C4004  ( .a(\prgm_register/en_not ), .b(a[307]), .out(
        \prgm_register/n616 ) );
  nand2 \prgm_register/C4005  ( .a(\prgm_register/n615 ), .b(
        \prgm_register/n616 ), .out(\prgm_register/or_signal [307]) );
  nand2 \prgm_register/C4006  ( .a(enable), .b(a[307]), .out(
        \prgm_register/n617 ) );
  nand2 \prgm_register/C4007  ( .a(\prgm_register/en_not ), .b(a[308]), .out(
        \prgm_register/n618 ) );
  nand2 \prgm_register/C4008  ( .a(\prgm_register/n617 ), .b(
        \prgm_register/n618 ), .out(\prgm_register/or_signal [308]) );
  nand2 \prgm_register/C4009  ( .a(enable), .b(a[308]), .out(
        \prgm_register/n619 ) );
  nand2 \prgm_register/C4010  ( .a(\prgm_register/en_not ), .b(a[309]), .out(
        \prgm_register/n620 ) );
  nand2 \prgm_register/C4011  ( .a(\prgm_register/n619 ), .b(
        \prgm_register/n620 ), .out(\prgm_register/or_signal [309]) );
  nand2 \prgm_register/C4012  ( .a(enable), .b(a[309]), .out(
        \prgm_register/n621 ) );
  nand2 \prgm_register/C4013  ( .a(\prgm_register/en_not ), .b(a[310]), .out(
        \prgm_register/n622 ) );
  nand2 \prgm_register/C4014  ( .a(\prgm_register/n621 ), .b(
        \prgm_register/n622 ), .out(\prgm_register/or_signal [310]) );
  nand2 \prgm_register/C4015  ( .a(enable), .b(a[310]), .out(
        \prgm_register/n623 ) );
  nand2 \prgm_register/C4016  ( .a(\prgm_register/en_not ), .b(a[311]), .out(
        \prgm_register/n624 ) );
  nand2 \prgm_register/C4017  ( .a(\prgm_register/n623 ), .b(
        \prgm_register/n624 ), .out(\prgm_register/or_signal [311]) );
  nand2 \prgm_register/C4018  ( .a(enable), .b(a[311]), .out(
        \prgm_register/n625 ) );
  nand2 \prgm_register/C4019  ( .a(\prgm_register/en_not ), .b(a[312]), .out(
        \prgm_register/n626 ) );
  nand2 \prgm_register/C4020  ( .a(\prgm_register/n625 ), .b(
        \prgm_register/n626 ), .out(\prgm_register/or_signal [312]) );
  nand2 \prgm_register/C4021  ( .a(enable), .b(a[312]), .out(
        \prgm_register/n627 ) );
  nand2 \prgm_register/C4022  ( .a(\prgm_register/en_not ), .b(a[313]), .out(
        \prgm_register/n628 ) );
  nand2 \prgm_register/C4023  ( .a(\prgm_register/n627 ), .b(
        \prgm_register/n628 ), .out(\prgm_register/or_signal [313]) );
  nand2 \prgm_register/C4024  ( .a(enable), .b(a[313]), .out(
        \prgm_register/n629 ) );
  nand2 \prgm_register/C4025  ( .a(\prgm_register/en_not ), .b(a[314]), .out(
        \prgm_register/n630 ) );
  nand2 \prgm_register/C4026  ( .a(\prgm_register/n629 ), .b(
        \prgm_register/n630 ), .out(\prgm_register/or_signal [314]) );
  nand2 \prgm_register/C4027  ( .a(enable), .b(a[314]), .out(
        \prgm_register/n631 ) );
  nand2 \prgm_register/C4028  ( .a(\prgm_register/en_not ), .b(a[315]), .out(
        \prgm_register/n632 ) );
  nand2 \prgm_register/C4029  ( .a(\prgm_register/n631 ), .b(
        \prgm_register/n632 ), .out(\prgm_register/or_signal [315]) );
  nand2 \prgm_register/C4030  ( .a(enable), .b(a[315]), .out(
        \prgm_register/n633 ) );
  nand2 \prgm_register/C4031  ( .a(\prgm_register/en_not ), .b(a[316]), .out(
        \prgm_register/n634 ) );
  nand2 \prgm_register/C4032  ( .a(\prgm_register/n633 ), .b(
        \prgm_register/n634 ), .out(\prgm_register/or_signal [316]) );
  nand2 \prgm_register/C4033  ( .a(enable), .b(a[316]), .out(
        \prgm_register/n635 ) );
  nand2 \prgm_register/C4034  ( .a(\prgm_register/en_not ), .b(a[317]), .out(
        \prgm_register/n636 ) );
  nand2 \prgm_register/C4035  ( .a(\prgm_register/n635 ), .b(
        \prgm_register/n636 ), .out(\prgm_register/or_signal [317]) );
  nand2 \prgm_register/C4036  ( .a(enable), .b(a[317]), .out(
        \prgm_register/n637 ) );
  nand2 \prgm_register/C4037  ( .a(\prgm_register/en_not ), .b(a[318]), .out(
        \prgm_register/n638 ) );
  nand2 \prgm_register/C4038  ( .a(\prgm_register/n637 ), .b(
        \prgm_register/n638 ), .out(\prgm_register/or_signal [318]) );
  nand2 \prgm_register/C4039  ( .a(enable), .b(a[318]), .out(
        \prgm_register/n639 ) );
  nand2 \prgm_register/C4040  ( .a(\prgm_register/en_not ), .b(a[319]), .out(
        \prgm_register/n640 ) );
  nand2 \prgm_register/C4041  ( .a(\prgm_register/n639 ), .b(
        \prgm_register/n640 ), .out(\prgm_register/or_signal [319]) );
  nand2 \prgm_register/C4042  ( .a(enable), .b(a[319]), .out(
        \prgm_register/n641 ) );
  nand2 \prgm_register/C4043  ( .a(\prgm_register/en_not ), .b(a[320]), .out(
        \prgm_register/n642 ) );
  nand2 \prgm_register/C4044  ( .a(\prgm_register/n641 ), .b(
        \prgm_register/n642 ), .out(\prgm_register/or_signal [320]) );
  nand2 \prgm_register/C4045  ( .a(enable), .b(a[320]), .out(
        \prgm_register/n643 ) );
  nand2 \prgm_register/C4046  ( .a(\prgm_register/en_not ), .b(a[321]), .out(
        \prgm_register/n644 ) );
  nand2 \prgm_register/C4047  ( .a(\prgm_register/n643 ), .b(
        \prgm_register/n644 ), .out(\prgm_register/or_signal [321]) );
  nand2 \prgm_register/C4048  ( .a(enable), .b(a[321]), .out(
        \prgm_register/n645 ) );
  nand2 \prgm_register/C4049  ( .a(\prgm_register/en_not ), .b(a[322]), .out(
        \prgm_register/n646 ) );
  nand2 \prgm_register/C4050  ( .a(\prgm_register/n645 ), .b(
        \prgm_register/n646 ), .out(\prgm_register/or_signal [322]) );
  nand2 \prgm_register/C4051  ( .a(enable), .b(a[322]), .out(
        \prgm_register/n647 ) );
  nand2 \prgm_register/C4052  ( .a(\prgm_register/en_not ), .b(a[323]), .out(
        \prgm_register/n648 ) );
  nand2 \prgm_register/C4053  ( .a(\prgm_register/n647 ), .b(
        \prgm_register/n648 ), .out(\prgm_register/or_signal [323]) );
  nand2 \prgm_register/C4054  ( .a(enable), .b(a[323]), .out(
        \prgm_register/n649 ) );
  nand2 \prgm_register/C4055  ( .a(\prgm_register/en_not ), .b(a[324]), .out(
        \prgm_register/n650 ) );
  nand2 \prgm_register/C4056  ( .a(\prgm_register/n649 ), .b(
        \prgm_register/n650 ), .out(\prgm_register/or_signal [324]) );
  nand2 \prgm_register/C4057  ( .a(enable), .b(a[324]), .out(
        \prgm_register/n651 ) );
  nand2 \prgm_register/C4058  ( .a(\prgm_register/en_not ), .b(a[325]), .out(
        \prgm_register/n652 ) );
  nand2 \prgm_register/C4059  ( .a(\prgm_register/n651 ), .b(
        \prgm_register/n652 ), .out(\prgm_register/or_signal [325]) );
  nand2 \prgm_register/C4060  ( .a(enable), .b(a[325]), .out(
        \prgm_register/n653 ) );
  nand2 \prgm_register/C4061  ( .a(\prgm_register/en_not ), .b(a[326]), .out(
        \prgm_register/n654 ) );
  nand2 \prgm_register/C4062  ( .a(\prgm_register/n653 ), .b(
        \prgm_register/n654 ), .out(\prgm_register/or_signal [326]) );
  nand2 \prgm_register/C4063  ( .a(enable), .b(a[326]), .out(
        \prgm_register/n655 ) );
  nand2 \prgm_register/C4064  ( .a(\prgm_register/en_not ), .b(a[327]), .out(
        \prgm_register/n656 ) );
  nand2 \prgm_register/C4065  ( .a(\prgm_register/n655 ), .b(
        \prgm_register/n656 ), .out(\prgm_register/or_signal [327]) );
  nand2 \prgm_register/C4066  ( .a(enable), .b(a[327]), .out(
        \prgm_register/n657 ) );
  nand2 \prgm_register/C4067  ( .a(\prgm_register/en_not ), .b(a[328]), .out(
        \prgm_register/n658 ) );
  nand2 \prgm_register/C4068  ( .a(\prgm_register/n657 ), .b(
        \prgm_register/n658 ), .out(\prgm_register/or_signal [328]) );
  nand2 \prgm_register/C4069  ( .a(enable), .b(a[328]), .out(
        \prgm_register/n659 ) );
  nand2 \prgm_register/C4070  ( .a(\prgm_register/en_not ), .b(a[329]), .out(
        \prgm_register/n660 ) );
  nand2 \prgm_register/C4071  ( .a(\prgm_register/n659 ), .b(
        \prgm_register/n660 ), .out(\prgm_register/or_signal [329]) );
  nand2 \prgm_register/C4072  ( .a(enable), .b(a[329]), .out(
        \prgm_register/n661 ) );
  nand2 \prgm_register/C4073  ( .a(\prgm_register/en_not ), .b(a[330]), .out(
        \prgm_register/n662 ) );
  nand2 \prgm_register/C4074  ( .a(\prgm_register/n661 ), .b(
        \prgm_register/n662 ), .out(\prgm_register/or_signal [330]) );
  nand2 \prgm_register/C4075  ( .a(enable), .b(a[330]), .out(
        \prgm_register/n663 ) );
  nand2 \prgm_register/C4076  ( .a(\prgm_register/en_not ), .b(a[331]), .out(
        \prgm_register/n664 ) );
  nand2 \prgm_register/C4077  ( .a(\prgm_register/n663 ), .b(
        \prgm_register/n664 ), .out(\prgm_register/or_signal [331]) );
  nand2 \prgm_register/C4078  ( .a(enable), .b(a[331]), .out(
        \prgm_register/n665 ) );
  nand2 \prgm_register/C4079  ( .a(\prgm_register/en_not ), .b(a[332]), .out(
        \prgm_register/n666 ) );
  nand2 \prgm_register/C4080  ( .a(\prgm_register/n665 ), .b(
        \prgm_register/n666 ), .out(\prgm_register/or_signal [332]) );
  nand2 \prgm_register/C4081  ( .a(enable), .b(a[332]), .out(
        \prgm_register/n667 ) );
  nand2 \prgm_register/C4082  ( .a(\prgm_register/en_not ), .b(a[333]), .out(
        \prgm_register/n668 ) );
  nand2 \prgm_register/C4083  ( .a(\prgm_register/n667 ), .b(
        \prgm_register/n668 ), .out(\prgm_register/or_signal [333]) );
  nand2 \prgm_register/C4084  ( .a(enable), .b(a[333]), .out(
        \prgm_register/n669 ) );
  nand2 \prgm_register/C4085  ( .a(\prgm_register/en_not ), .b(a[334]), .out(
        \prgm_register/n670 ) );
  nand2 \prgm_register/C4086  ( .a(\prgm_register/n669 ), .b(
        \prgm_register/n670 ), .out(\prgm_register/or_signal [334]) );
  nand2 \prgm_register/C4087  ( .a(enable), .b(a[334]), .out(
        \prgm_register/n671 ) );
  nand2 \prgm_register/C4088  ( .a(\prgm_register/en_not ), .b(a[335]), .out(
        \prgm_register/n672 ) );
  nand2 \prgm_register/C4089  ( .a(\prgm_register/n671 ), .b(
        \prgm_register/n672 ), .out(\prgm_register/or_signal [335]) );
  nand2 \prgm_register/C4090  ( .a(enable), .b(a[335]), .out(
        \prgm_register/n673 ) );
  nand2 \prgm_register/C4091  ( .a(\prgm_register/en_not ), .b(a[336]), .out(
        \prgm_register/n674 ) );
  nand2 \prgm_register/C4092  ( .a(\prgm_register/n673 ), .b(
        \prgm_register/n674 ), .out(\prgm_register/or_signal [336]) );
  nand2 \prgm_register/C4093  ( .a(enable), .b(a[336]), .out(
        \prgm_register/n675 ) );
  nand2 \prgm_register/C4094  ( .a(\prgm_register/en_not ), .b(a[337]), .out(
        \prgm_register/n676 ) );
  nand2 \prgm_register/C4095  ( .a(\prgm_register/n675 ), .b(
        \prgm_register/n676 ), .out(\prgm_register/or_signal [337]) );
  nand2 \prgm_register/C4096  ( .a(enable), .b(a[337]), .out(
        \prgm_register/n677 ) );
  nand2 \prgm_register/C4097  ( .a(\prgm_register/en_not ), .b(a[338]), .out(
        \prgm_register/n678 ) );
  nand2 \prgm_register/C4098  ( .a(\prgm_register/n677 ), .b(
        \prgm_register/n678 ), .out(\prgm_register/or_signal [338]) );
  nand2 \prgm_register/C4099  ( .a(enable), .b(a[338]), .out(
        \prgm_register/n679 ) );
  nand2 \prgm_register/C4100  ( .a(\prgm_register/en_not ), .b(a[339]), .out(
        \prgm_register/n680 ) );
  nand2 \prgm_register/C4101  ( .a(\prgm_register/n679 ), .b(
        \prgm_register/n680 ), .out(\prgm_register/or_signal [339]) );
  nand2 \prgm_register/C4102  ( .a(enable), .b(a[339]), .out(
        \prgm_register/n681 ) );
  nand2 \prgm_register/C4103  ( .a(\prgm_register/en_not ), .b(a[340]), .out(
        \prgm_register/n682 ) );
  nand2 \prgm_register/C4104  ( .a(\prgm_register/n681 ), .b(
        \prgm_register/n682 ), .out(\prgm_register/or_signal [340]) );
  nand2 \prgm_register/C4105  ( .a(enable), .b(a[340]), .out(
        \prgm_register/n683 ) );
  nand2 \prgm_register/C4106  ( .a(\prgm_register/en_not ), .b(a[341]), .out(
        \prgm_register/n684 ) );
  nand2 \prgm_register/C4107  ( .a(\prgm_register/n683 ), .b(
        \prgm_register/n684 ), .out(\prgm_register/or_signal [341]) );
  nand2 \prgm_register/C4108  ( .a(enable), .b(a[341]), .out(
        \prgm_register/n685 ) );
  nand2 \prgm_register/C4109  ( .a(\prgm_register/en_not ), .b(a[342]), .out(
        \prgm_register/n686 ) );
  nand2 \prgm_register/C4110  ( .a(\prgm_register/n685 ), .b(
        \prgm_register/n686 ), .out(\prgm_register/or_signal [342]) );
  nand2 \prgm_register/C4111  ( .a(enable), .b(a[342]), .out(
        \prgm_register/n687 ) );
  nand2 \prgm_register/C4112  ( .a(\prgm_register/en_not ), .b(a[343]), .out(
        \prgm_register/n688 ) );
  nand2 \prgm_register/C4113  ( .a(\prgm_register/n687 ), .b(
        \prgm_register/n688 ), .out(\prgm_register/or_signal [343]) );
  nand2 \prgm_register/C4114  ( .a(enable), .b(a[343]), .out(
        \prgm_register/n689 ) );
  nand2 \prgm_register/C4115  ( .a(\prgm_register/en_not ), .b(a[344]), .out(
        \prgm_register/n690 ) );
  nand2 \prgm_register/C4116  ( .a(\prgm_register/n689 ), .b(
        \prgm_register/n690 ), .out(\prgm_register/or_signal [344]) );
  nand2 \prgm_register/C4117  ( .a(enable), .b(a[344]), .out(
        \prgm_register/n691 ) );
  nand2 \prgm_register/C4118  ( .a(\prgm_register/en_not ), .b(a[345]), .out(
        \prgm_register/n692 ) );
  nand2 \prgm_register/C4119  ( .a(\prgm_register/n691 ), .b(
        \prgm_register/n692 ), .out(\prgm_register/or_signal [345]) );
  nand2 \prgm_register/C4120  ( .a(enable), .b(a[345]), .out(
        \prgm_register/n693 ) );
  nand2 \prgm_register/C4121  ( .a(\prgm_register/en_not ), .b(a[346]), .out(
        \prgm_register/n694 ) );
  nand2 \prgm_register/C4122  ( .a(\prgm_register/n693 ), .b(
        \prgm_register/n694 ), .out(\prgm_register/or_signal [346]) );
  nand2 \prgm_register/C4123  ( .a(enable), .b(a[346]), .out(
        \prgm_register/n695 ) );
  nand2 \prgm_register/C4124  ( .a(\prgm_register/en_not ), .b(a[347]), .out(
        \prgm_register/n696 ) );
  nand2 \prgm_register/C4125  ( .a(\prgm_register/n695 ), .b(
        \prgm_register/n696 ), .out(\prgm_register/or_signal [347]) );
  nand2 \prgm_register/C4126  ( .a(enable), .b(a[347]), .out(
        \prgm_register/n697 ) );
  nand2 \prgm_register/C4127  ( .a(\prgm_register/en_not ), .b(a[348]), .out(
        \prgm_register/n698 ) );
  nand2 \prgm_register/C4128  ( .a(\prgm_register/n697 ), .b(
        \prgm_register/n698 ), .out(\prgm_register/or_signal [348]) );
  nand2 \prgm_register/C4129  ( .a(enable), .b(a[348]), .out(
        \prgm_register/n699 ) );
  nand2 \prgm_register/C4130  ( .a(\prgm_register/en_not ), .b(a[349]), .out(
        \prgm_register/n700 ) );
  nand2 \prgm_register/C4131  ( .a(\prgm_register/n699 ), .b(
        \prgm_register/n700 ), .out(\prgm_register/or_signal [349]) );
  nand2 \prgm_register/C4132  ( .a(enable), .b(a[349]), .out(
        \prgm_register/n701 ) );
  nand2 \prgm_register/C4133  ( .a(\prgm_register/en_not ), .b(a[350]), .out(
        \prgm_register/n702 ) );
  nand2 \prgm_register/C4134  ( .a(\prgm_register/n701 ), .b(
        \prgm_register/n702 ), .out(\prgm_register/or_signal [350]) );
  nand2 \prgm_register/C4135  ( .a(enable), .b(a[350]), .out(
        \prgm_register/n703 ) );
  nand2 \prgm_register/C4136  ( .a(\prgm_register/en_not ), .b(a[351]), .out(
        \prgm_register/n704 ) );
  nand2 \prgm_register/C4137  ( .a(\prgm_register/n703 ), .b(
        \prgm_register/n704 ), .out(\prgm_register/or_signal [351]) );
  nand2 \prgm_register/C4138  ( .a(enable), .b(a[351]), .out(
        \prgm_register/n705 ) );
  nand2 \prgm_register/C4139  ( .a(\prgm_register/en_not ), .b(a[352]), .out(
        \prgm_register/n706 ) );
  nand2 \prgm_register/C4140  ( .a(\prgm_register/n705 ), .b(
        \prgm_register/n706 ), .out(\prgm_register/or_signal [352]) );
  nand2 \prgm_register/C4141  ( .a(enable), .b(a[352]), .out(
        \prgm_register/n707 ) );
  nand2 \prgm_register/C4142  ( .a(\prgm_register/en_not ), .b(a[353]), .out(
        \prgm_register/n708 ) );
  nand2 \prgm_register/C4143  ( .a(\prgm_register/n707 ), .b(
        \prgm_register/n708 ), .out(\prgm_register/or_signal [353]) );
  nand2 \prgm_register/C4144  ( .a(enable), .b(a[353]), .out(
        \prgm_register/n709 ) );
  nand2 \prgm_register/C4145  ( .a(\prgm_register/en_not ), .b(a[354]), .out(
        \prgm_register/n710 ) );
  nand2 \prgm_register/C4146  ( .a(\prgm_register/n709 ), .b(
        \prgm_register/n710 ), .out(\prgm_register/or_signal [354]) );
  nand2 \prgm_register/C4147  ( .a(enable), .b(a[354]), .out(
        \prgm_register/n711 ) );
  nand2 \prgm_register/C4148  ( .a(\prgm_register/en_not ), .b(a[355]), .out(
        \prgm_register/n712 ) );
  nand2 \prgm_register/C4149  ( .a(\prgm_register/n711 ), .b(
        \prgm_register/n712 ), .out(\prgm_register/or_signal [355]) );
  nand2 \prgm_register/C4150  ( .a(enable), .b(a[355]), .out(
        \prgm_register/n713 ) );
  nand2 \prgm_register/C4151  ( .a(\prgm_register/en_not ), .b(a[356]), .out(
        \prgm_register/n714 ) );
  nand2 \prgm_register/C4152  ( .a(\prgm_register/n713 ), .b(
        \prgm_register/n714 ), .out(\prgm_register/or_signal [356]) );
  nand2 \prgm_register/C4153  ( .a(enable), .b(a[356]), .out(
        \prgm_register/n715 ) );
  nand2 \prgm_register/C4154  ( .a(\prgm_register/en_not ), .b(a[357]), .out(
        \prgm_register/n716 ) );
  nand2 \prgm_register/C4155  ( .a(\prgm_register/n715 ), .b(
        \prgm_register/n716 ), .out(\prgm_register/or_signal [357]) );
  nand2 \prgm_register/C4156  ( .a(enable), .b(a[357]), .out(
        \prgm_register/n717 ) );
  nand2 \prgm_register/C4157  ( .a(\prgm_register/en_not ), .b(a[358]), .out(
        \prgm_register/n718 ) );
  nand2 \prgm_register/C4158  ( .a(\prgm_register/n717 ), .b(
        \prgm_register/n718 ), .out(\prgm_register/or_signal [358]) );
  nand2 \prgm_register/C4159  ( .a(enable), .b(a[358]), .out(
        \prgm_register/n719 ) );
  nand2 \prgm_register/C4160  ( .a(\prgm_register/en_not ), .b(a[359]), .out(
        \prgm_register/n720 ) );
  nand2 \prgm_register/C4161  ( .a(\prgm_register/n719 ), .b(
        \prgm_register/n720 ), .out(\prgm_register/or_signal [359]) );
  nand2 \prgm_register/C4162  ( .a(enable), .b(a[359]), .out(
        \prgm_register/n721 ) );
  nand2 \prgm_register/C4163  ( .a(\prgm_register/en_not ), .b(a[360]), .out(
        \prgm_register/n722 ) );
  nand2 \prgm_register/C4164  ( .a(\prgm_register/n721 ), .b(
        \prgm_register/n722 ), .out(\prgm_register/or_signal [360]) );
  nand2 \prgm_register/C4165  ( .a(enable), .b(a[360]), .out(
        \prgm_register/n723 ) );
  nand2 \prgm_register/C4166  ( .a(\prgm_register/en_not ), .b(a[361]), .out(
        \prgm_register/n724 ) );
  nand2 \prgm_register/C4167  ( .a(\prgm_register/n723 ), .b(
        \prgm_register/n724 ), .out(\prgm_register/or_signal [361]) );
  nand2 \prgm_register/C4168  ( .a(enable), .b(a[361]), .out(
        \prgm_register/n725 ) );
  nand2 \prgm_register/C4169  ( .a(\prgm_register/en_not ), .b(a[362]), .out(
        \prgm_register/n726 ) );
  nand2 \prgm_register/C4170  ( .a(\prgm_register/n725 ), .b(
        \prgm_register/n726 ), .out(\prgm_register/or_signal [362]) );
  nand2 \prgm_register/C4171  ( .a(enable), .b(a[362]), .out(
        \prgm_register/n727 ) );
  nand2 \prgm_register/C4172  ( .a(\prgm_register/en_not ), .b(a[363]), .out(
        \prgm_register/n728 ) );
  nand2 \prgm_register/C4173  ( .a(\prgm_register/n727 ), .b(
        \prgm_register/n728 ), .out(\prgm_register/or_signal [363]) );
  nand2 \prgm_register/C4174  ( .a(enable), .b(a[363]), .out(
        \prgm_register/n729 ) );
  nand2 \prgm_register/C4175  ( .a(\prgm_register/en_not ), .b(a[364]), .out(
        \prgm_register/n730 ) );
  nand2 \prgm_register/C4176  ( .a(\prgm_register/n729 ), .b(
        \prgm_register/n730 ), .out(\prgm_register/or_signal [364]) );
  nand2 \prgm_register/C4177  ( .a(enable), .b(a[364]), .out(
        \prgm_register/n731 ) );
  nand2 \prgm_register/C4178  ( .a(\prgm_register/en_not ), .b(a[365]), .out(
        \prgm_register/n732 ) );
  nand2 \prgm_register/C4179  ( .a(\prgm_register/n731 ), .b(
        \prgm_register/n732 ), .out(\prgm_register/or_signal [365]) );
  nand2 \prgm_register/C4180  ( .a(enable), .b(a[365]), .out(
        \prgm_register/n733 ) );
  nand2 \prgm_register/C4181  ( .a(\prgm_register/en_not ), .b(a[366]), .out(
        \prgm_register/n734 ) );
  nand2 \prgm_register/C4182  ( .a(\prgm_register/n733 ), .b(
        \prgm_register/n734 ), .out(\prgm_register/or_signal [366]) );
  nand2 \prgm_register/C4183  ( .a(enable), .b(a[366]), .out(
        \prgm_register/n735 ) );
  nand2 \prgm_register/C4184  ( .a(\prgm_register/en_not ), .b(a[367]), .out(
        \prgm_register/n736 ) );
  nand2 \prgm_register/C4185  ( .a(\prgm_register/n735 ), .b(
        \prgm_register/n736 ), .out(\prgm_register/or_signal [367]) );
  nand2 \prgm_register/C4186  ( .a(enable), .b(a[367]), .out(
        \prgm_register/n737 ) );
  nand2 \prgm_register/C4187  ( .a(\prgm_register/en_not ), .b(a[368]), .out(
        \prgm_register/n738 ) );
  nand2 \prgm_register/C4188  ( .a(\prgm_register/n737 ), .b(
        \prgm_register/n738 ), .out(\prgm_register/or_signal [368]) );
  nand2 \prgm_register/C4189  ( .a(enable), .b(a[368]), .out(
        \prgm_register/n739 ) );
  nand2 \prgm_register/C4190  ( .a(\prgm_register/en_not ), .b(a[369]), .out(
        \prgm_register/n740 ) );
  nand2 \prgm_register/C4191  ( .a(\prgm_register/n739 ), .b(
        \prgm_register/n740 ), .out(\prgm_register/or_signal [369]) );
  nand2 \prgm_register/C4192  ( .a(enable), .b(a[369]), .out(
        \prgm_register/n741 ) );
  nand2 \prgm_register/C4193  ( .a(\prgm_register/en_not ), .b(a[370]), .out(
        \prgm_register/n742 ) );
  nand2 \prgm_register/C4194  ( .a(\prgm_register/n741 ), .b(
        \prgm_register/n742 ), .out(\prgm_register/or_signal [370]) );
  nand2 \prgm_register/C4195  ( .a(enable), .b(a[370]), .out(
        \prgm_register/n743 ) );
  nand2 \prgm_register/C4196  ( .a(\prgm_register/en_not ), .b(a[371]), .out(
        \prgm_register/n744 ) );
  nand2 \prgm_register/C4197  ( .a(\prgm_register/n743 ), .b(
        \prgm_register/n744 ), .out(\prgm_register/or_signal [371]) );
  nand2 \prgm_register/C4198  ( .a(enable), .b(a[371]), .out(
        \prgm_register/n745 ) );
  nand2 \prgm_register/C4199  ( .a(\prgm_register/en_not ), .b(a[372]), .out(
        \prgm_register/n746 ) );
  nand2 \prgm_register/C4200  ( .a(\prgm_register/n745 ), .b(
        \prgm_register/n746 ), .out(\prgm_register/or_signal [372]) );
  nand2 \prgm_register/C4201  ( .a(enable), .b(a[372]), .out(
        \prgm_register/n747 ) );
  nand2 \prgm_register/C4202  ( .a(\prgm_register/en_not ), .b(a[373]), .out(
        \prgm_register/n748 ) );
  nand2 \prgm_register/C4203  ( .a(\prgm_register/n747 ), .b(
        \prgm_register/n748 ), .out(\prgm_register/or_signal [373]) );
  nand2 \prgm_register/C4204  ( .a(enable), .b(a[373]), .out(
        \prgm_register/n749 ) );
  nand2 \prgm_register/C4205  ( .a(\prgm_register/en_not ), .b(a[374]), .out(
        \prgm_register/n750 ) );
  nand2 \prgm_register/C4206  ( .a(\prgm_register/n749 ), .b(
        \prgm_register/n750 ), .out(\prgm_register/or_signal [374]) );
  nand2 \prgm_register/C4207  ( .a(enable), .b(a[374]), .out(
        \prgm_register/n751 ) );
  nand2 \prgm_register/C4208  ( .a(\prgm_register/en_not ), .b(a[375]), .out(
        \prgm_register/n752 ) );
  nand2 \prgm_register/C4209  ( .a(\prgm_register/n751 ), .b(
        \prgm_register/n752 ), .out(\prgm_register/or_signal [375]) );
  nand2 \prgm_register/C4210  ( .a(enable), .b(a[375]), .out(
        \prgm_register/n753 ) );
  nand2 \prgm_register/C4211  ( .a(\prgm_register/en_not ), .b(a[376]), .out(
        \prgm_register/n754 ) );
  nand2 \prgm_register/C4212  ( .a(\prgm_register/n753 ), .b(
        \prgm_register/n754 ), .out(\prgm_register/or_signal [376]) );
  nand2 \prgm_register/C4213  ( .a(enable), .b(a[376]), .out(
        \prgm_register/n755 ) );
  nand2 \prgm_register/C4214  ( .a(\prgm_register/en_not ), .b(a[377]), .out(
        \prgm_register/n756 ) );
  nand2 \prgm_register/C4215  ( .a(\prgm_register/n755 ), .b(
        \prgm_register/n756 ), .out(\prgm_register/or_signal [377]) );
  nand2 \prgm_register/C4216  ( .a(enable), .b(a[377]), .out(
        \prgm_register/n757 ) );
  nand2 \prgm_register/C4217  ( .a(\prgm_register/en_not ), .b(a[378]), .out(
        \prgm_register/n758 ) );
  nand2 \prgm_register/C4218  ( .a(\prgm_register/n757 ), .b(
        \prgm_register/n758 ), .out(\prgm_register/or_signal [378]) );
  nand2 \prgm_register/C4219  ( .a(enable), .b(a[378]), .out(
        \prgm_register/n759 ) );
  nand2 \prgm_register/C4220  ( .a(\prgm_register/en_not ), .b(a[379]), .out(
        \prgm_register/n760 ) );
  nand2 \prgm_register/C4221  ( .a(\prgm_register/n759 ), .b(
        \prgm_register/n760 ), .out(\prgm_register/or_signal [379]) );
  nand2 \prgm_register/C4222  ( .a(enable), .b(a[379]), .out(
        \prgm_register/n761 ) );
  nand2 \prgm_register/C4223  ( .a(\prgm_register/en_not ), .b(a[380]), .out(
        \prgm_register/n762 ) );
  nand2 \prgm_register/C4224  ( .a(\prgm_register/n761 ), .b(
        \prgm_register/n762 ), .out(\prgm_register/or_signal [380]) );
  nand2 \prgm_register/C4225  ( .a(enable), .b(a[380]), .out(
        \prgm_register/n763 ) );
  nand2 \prgm_register/C4226  ( .a(\prgm_register/en_not ), .b(a[381]), .out(
        \prgm_register/n764 ) );
  nand2 \prgm_register/C4227  ( .a(\prgm_register/n763 ), .b(
        \prgm_register/n764 ), .out(\prgm_register/or_signal [381]) );
  nand2 \prgm_register/C4228  ( .a(enable), .b(a[381]), .out(
        \prgm_register/n765 ) );
  nand2 \prgm_register/C4229  ( .a(\prgm_register/en_not ), .b(a[382]), .out(
        \prgm_register/n766 ) );
  nand2 \prgm_register/C4230  ( .a(\prgm_register/n765 ), .b(
        \prgm_register/n766 ), .out(\prgm_register/or_signal [382]) );
  nand2 \prgm_register/C4231  ( .a(enable), .b(a[382]), .out(
        \prgm_register/n767 ) );
  nand2 \prgm_register/C4232  ( .a(\prgm_register/en_not ), .b(a[383]), .out(
        \prgm_register/n768 ) );
  nand2 \prgm_register/C4233  ( .a(\prgm_register/n767 ), .b(
        \prgm_register/n768 ), .out(\prgm_register/or_signal [383]) );
  nand2 \prgm_register/C4234  ( .a(enable), .b(a[383]), .out(
        \prgm_register/n769 ) );
  nand2 \prgm_register/C4235  ( .a(\prgm_register/en_not ), .b(a[384]), .out(
        \prgm_register/n770 ) );
  nand2 \prgm_register/C4236  ( .a(\prgm_register/n769 ), .b(
        \prgm_register/n770 ), .out(\prgm_register/or_signal [384]) );
  nand2 \prgm_register/C4237  ( .a(enable), .b(a[384]), .out(
        \prgm_register/n771 ) );
  nand2 \prgm_register/C4238  ( .a(\prgm_register/en_not ), .b(a[385]), .out(
        \prgm_register/n772 ) );
  nand2 \prgm_register/C4239  ( .a(\prgm_register/n771 ), .b(
        \prgm_register/n772 ), .out(\prgm_register/or_signal [385]) );
  nand2 \prgm_register/C4240  ( .a(enable), .b(a[385]), .out(
        \prgm_register/n773 ) );
  nand2 \prgm_register/C4241  ( .a(\prgm_register/en_not ), .b(a[386]), .out(
        \prgm_register/n774 ) );
  nand2 \prgm_register/C4242  ( .a(\prgm_register/n773 ), .b(
        \prgm_register/n774 ), .out(\prgm_register/or_signal [386]) );
  nand2 \prgm_register/C4243  ( .a(enable), .b(a[386]), .out(
        \prgm_register/n775 ) );
  nand2 \prgm_register/C4244  ( .a(\prgm_register/en_not ), .b(a[387]), .out(
        \prgm_register/n776 ) );
  nand2 \prgm_register/C4245  ( .a(\prgm_register/n775 ), .b(
        \prgm_register/n776 ), .out(\prgm_register/or_signal [387]) );
  nand2 \prgm_register/C4246  ( .a(enable), .b(a[387]), .out(
        \prgm_register/n777 ) );
  nand2 \prgm_register/C4247  ( .a(\prgm_register/en_not ), .b(a[388]), .out(
        \prgm_register/n778 ) );
  nand2 \prgm_register/C4248  ( .a(\prgm_register/n777 ), .b(
        \prgm_register/n778 ), .out(\prgm_register/or_signal [388]) );
  nand2 \prgm_register/C4249  ( .a(enable), .b(a[388]), .out(
        \prgm_register/n779 ) );
  nand2 \prgm_register/C4250  ( .a(\prgm_register/en_not ), .b(a[389]), .out(
        \prgm_register/n780 ) );
  nand2 \prgm_register/C4251  ( .a(\prgm_register/n779 ), .b(
        \prgm_register/n780 ), .out(\prgm_register/or_signal [389]) );
  nand2 \prgm_register/C4252  ( .a(enable), .b(a[389]), .out(
        \prgm_register/n781 ) );
  nand2 \prgm_register/C4253  ( .a(\prgm_register/en_not ), .b(a[390]), .out(
        \prgm_register/n782 ) );
  nand2 \prgm_register/C4254  ( .a(\prgm_register/n781 ), .b(
        \prgm_register/n782 ), .out(\prgm_register/or_signal [390]) );
  nand2 \prgm_register/C4255  ( .a(enable), .b(a[390]), .out(
        \prgm_register/n783 ) );
  nand2 \prgm_register/C4256  ( .a(\prgm_register/en_not ), .b(a[391]), .out(
        \prgm_register/n784 ) );
  nand2 \prgm_register/C4257  ( .a(\prgm_register/n783 ), .b(
        \prgm_register/n784 ), .out(\prgm_register/or_signal [391]) );
  nand2 \prgm_register/C4258  ( .a(enable), .b(a[391]), .out(
        \prgm_register/n785 ) );
  nand2 \prgm_register/C4259  ( .a(\prgm_register/en_not ), .b(a[392]), .out(
        \prgm_register/n786 ) );
  nand2 \prgm_register/C4260  ( .a(\prgm_register/n785 ), .b(
        \prgm_register/n786 ), .out(\prgm_register/or_signal [392]) );
  nand2 \prgm_register/C4261  ( .a(enable), .b(a[392]), .out(
        \prgm_register/n787 ) );
  nand2 \prgm_register/C4262  ( .a(\prgm_register/en_not ), .b(a[393]), .out(
        \prgm_register/n788 ) );
  nand2 \prgm_register/C4263  ( .a(\prgm_register/n787 ), .b(
        \prgm_register/n788 ), .out(\prgm_register/or_signal [393]) );
  nand2 \prgm_register/C4264  ( .a(enable), .b(a[393]), .out(
        \prgm_register/n789 ) );
  nand2 \prgm_register/C4265  ( .a(\prgm_register/en_not ), .b(a[394]), .out(
        \prgm_register/n790 ) );
  nand2 \prgm_register/C4266  ( .a(\prgm_register/n789 ), .b(
        \prgm_register/n790 ), .out(\prgm_register/or_signal [394]) );
  nand2 \prgm_register/C4267  ( .a(enable), .b(a[394]), .out(
        \prgm_register/n791 ) );
  nand2 \prgm_register/C4268  ( .a(\prgm_register/en_not ), .b(a[395]), .out(
        \prgm_register/n792 ) );
  nand2 \prgm_register/C4269  ( .a(\prgm_register/n791 ), .b(
        \prgm_register/n792 ), .out(\prgm_register/or_signal [395]) );
  nand2 \prgm_register/C4270  ( .a(enable), .b(a[395]), .out(
        \prgm_register/n793 ) );
  nand2 \prgm_register/C4271  ( .a(\prgm_register/en_not ), .b(a[396]), .out(
        \prgm_register/n794 ) );
  nand2 \prgm_register/C4272  ( .a(\prgm_register/n793 ), .b(
        \prgm_register/n794 ), .out(\prgm_register/or_signal [396]) );
  nand2 \prgm_register/C4273  ( .a(enable), .b(a[396]), .out(
        \prgm_register/n795 ) );
  nand2 \prgm_register/C4274  ( .a(\prgm_register/en_not ), .b(a[397]), .out(
        \prgm_register/n796 ) );
  nand2 \prgm_register/C4275  ( .a(\prgm_register/n795 ), .b(
        \prgm_register/n796 ), .out(\prgm_register/or_signal [397]) );
  nand2 \prgm_register/C4276  ( .a(enable), .b(a[397]), .out(
        \prgm_register/n797 ) );
  nand2 \prgm_register/C4277  ( .a(\prgm_register/en_not ), .b(a[398]), .out(
        \prgm_register/n798 ) );
  nand2 \prgm_register/C4278  ( .a(\prgm_register/n797 ), .b(
        \prgm_register/n798 ), .out(\prgm_register/or_signal [398]) );
  nand2 \prgm_register/C4279  ( .a(enable), .b(a[398]), .out(
        \prgm_register/n799 ) );
  nand2 \prgm_register/C4280  ( .a(\prgm_register/en_not ), .b(a[399]), .out(
        \prgm_register/n800 ) );
  nand2 \prgm_register/C4281  ( .a(\prgm_register/n799 ), .b(
        \prgm_register/n800 ), .out(\prgm_register/or_signal [399]) );
  nand2 \prgm_register/C4282  ( .a(enable), .b(a[399]), .out(
        \prgm_register/n801 ) );
  nand2 \prgm_register/C4283  ( .a(\prgm_register/en_not ), .b(a[400]), .out(
        \prgm_register/n802 ) );
  nand2 \prgm_register/C4284  ( .a(\prgm_register/n801 ), .b(
        \prgm_register/n802 ), .out(\prgm_register/or_signal [400]) );
  nand2 \prgm_register/C4285  ( .a(enable), .b(a[400]), .out(
        \prgm_register/n803 ) );
  nand2 \prgm_register/C4286  ( .a(\prgm_register/en_not ), .b(a[401]), .out(
        \prgm_register/n804 ) );
  nand2 \prgm_register/C4287  ( .a(\prgm_register/n803 ), .b(
        \prgm_register/n804 ), .out(\prgm_register/or_signal [401]) );
  nand2 \prgm_register/C4288  ( .a(enable), .b(a[401]), .out(
        \prgm_register/n805 ) );
  nand2 \prgm_register/C4289  ( .a(\prgm_register/en_not ), .b(a[402]), .out(
        \prgm_register/n806 ) );
  nand2 \prgm_register/C4290  ( .a(\prgm_register/n805 ), .b(
        \prgm_register/n806 ), .out(\prgm_register/or_signal [402]) );
  nand2 \prgm_register/C4291  ( .a(enable), .b(a[402]), .out(
        \prgm_register/n807 ) );
  nand2 \prgm_register/C4292  ( .a(\prgm_register/en_not ), .b(a[403]), .out(
        \prgm_register/n808 ) );
  nand2 \prgm_register/C4293  ( .a(\prgm_register/n807 ), .b(
        \prgm_register/n808 ), .out(\prgm_register/or_signal [403]) );
  nand2 \prgm_register/C4294  ( .a(enable), .b(a[403]), .out(
        \prgm_register/n809 ) );
  nand2 \prgm_register/C4295  ( .a(\prgm_register/en_not ), .b(a[404]), .out(
        \prgm_register/n810 ) );
  nand2 \prgm_register/C4296  ( .a(\prgm_register/n809 ), .b(
        \prgm_register/n810 ), .out(\prgm_register/or_signal [404]) );
  nand2 \prgm_register/C4297  ( .a(enable), .b(a[404]), .out(
        \prgm_register/n811 ) );
  nand2 \prgm_register/C4298  ( .a(\prgm_register/en_not ), .b(a[405]), .out(
        \prgm_register/n812 ) );
  nand2 \prgm_register/C4299  ( .a(\prgm_register/n811 ), .b(
        \prgm_register/n812 ), .out(\prgm_register/or_signal [405]) );
  nand2 \prgm_register/C4300  ( .a(enable), .b(a[405]), .out(
        \prgm_register/n813 ) );
  nand2 \prgm_register/C4301  ( .a(\prgm_register/en_not ), .b(a[406]), .out(
        \prgm_register/n814 ) );
  nand2 \prgm_register/C4302  ( .a(\prgm_register/n813 ), .b(
        \prgm_register/n814 ), .out(\prgm_register/or_signal [406]) );
  nand2 \prgm_register/C4303  ( .a(enable), .b(a[406]), .out(
        \prgm_register/n815 ) );
  nand2 \prgm_register/C4304  ( .a(\prgm_register/en_not ), .b(a[407]), .out(
        \prgm_register/n816 ) );
  nand2 \prgm_register/C4305  ( .a(\prgm_register/n815 ), .b(
        \prgm_register/n816 ), .out(\prgm_register/or_signal [407]) );
  nand2 \prgm_register/C4306  ( .a(enable), .b(a[407]), .out(
        \prgm_register/n817 ) );
  nand2 \prgm_register/C4307  ( .a(\prgm_register/en_not ), .b(a[408]), .out(
        \prgm_register/n818 ) );
  nand2 \prgm_register/C4308  ( .a(\prgm_register/n817 ), .b(
        \prgm_register/n818 ), .out(\prgm_register/or_signal [408]) );
  nand2 \prgm_register/C4309  ( .a(enable), .b(a[408]), .out(
        \prgm_register/n819 ) );
  nand2 \prgm_register/C4310  ( .a(\prgm_register/en_not ), .b(a[409]), .out(
        \prgm_register/n820 ) );
  nand2 \prgm_register/C4311  ( .a(\prgm_register/n819 ), .b(
        \prgm_register/n820 ), .out(\prgm_register/or_signal [409]) );
  nand2 \prgm_register/C4312  ( .a(enable), .b(a[409]), .out(
        \prgm_register/n821 ) );
  nand2 \prgm_register/C4313  ( .a(\prgm_register/en_not ), .b(a[410]), .out(
        \prgm_register/n822 ) );
  nand2 \prgm_register/C4314  ( .a(\prgm_register/n821 ), .b(
        \prgm_register/n822 ), .out(\prgm_register/or_signal [410]) );
  nand2 \prgm_register/C4315  ( .a(enable), .b(a[410]), .out(
        \prgm_register/n823 ) );
  nand2 \prgm_register/C4316  ( .a(\prgm_register/en_not ), .b(a[411]), .out(
        \prgm_register/n824 ) );
  nand2 \prgm_register/C4317  ( .a(\prgm_register/n823 ), .b(
        \prgm_register/n824 ), .out(\prgm_register/or_signal [411]) );
  nand2 \prgm_register/C4318  ( .a(enable), .b(a[411]), .out(
        \prgm_register/n825 ) );
  nand2 \prgm_register/C4319  ( .a(\prgm_register/en_not ), .b(a[412]), .out(
        \prgm_register/n826 ) );
  nand2 \prgm_register/C4320  ( .a(\prgm_register/n825 ), .b(
        \prgm_register/n826 ), .out(\prgm_register/or_signal [412]) );
  nand2 \prgm_register/C4321  ( .a(enable), .b(a[412]), .out(
        \prgm_register/n827 ) );
  nand2 \prgm_register/C4322  ( .a(\prgm_register/en_not ), .b(a[413]), .out(
        \prgm_register/n828 ) );
  nand2 \prgm_register/C4323  ( .a(\prgm_register/n827 ), .b(
        \prgm_register/n828 ), .out(\prgm_register/or_signal [413]) );
  nand2 \prgm_register/C4324  ( .a(enable), .b(a[413]), .out(
        \prgm_register/n829 ) );
  nand2 \prgm_register/C4325  ( .a(\prgm_register/en_not ), .b(a[414]), .out(
        \prgm_register/n830 ) );
  nand2 \prgm_register/C4326  ( .a(\prgm_register/n829 ), .b(
        \prgm_register/n830 ), .out(\prgm_register/or_signal [414]) );
  nand2 \prgm_register/C4327  ( .a(enable), .b(a[414]), .out(
        \prgm_register/n831 ) );
  nand2 \prgm_register/C4328  ( .a(\prgm_register/en_not ), .b(a[415]), .out(
        \prgm_register/n832 ) );
  nand2 \prgm_register/C4329  ( .a(\prgm_register/n831 ), .b(
        \prgm_register/n832 ), .out(\prgm_register/or_signal [415]) );
  nand2 \prgm_register/C4330  ( .a(enable), .b(a[415]), .out(
        \prgm_register/n833 ) );
  nand2 \prgm_register/C4331  ( .a(\prgm_register/en_not ), .b(a[416]), .out(
        \prgm_register/n834 ) );
  nand2 \prgm_register/C4332  ( .a(\prgm_register/n833 ), .b(
        \prgm_register/n834 ), .out(\prgm_register/or_signal [416]) );
  nand2 \prgm_register/C4333  ( .a(enable), .b(a[416]), .out(
        \prgm_register/n835 ) );
  nand2 \prgm_register/C4334  ( .a(\prgm_register/en_not ), .b(a[417]), .out(
        \prgm_register/n836 ) );
  nand2 \prgm_register/C4335  ( .a(\prgm_register/n835 ), .b(
        \prgm_register/n836 ), .out(\prgm_register/or_signal [417]) );
  nand2 \prgm_register/C4336  ( .a(enable), .b(a[417]), .out(
        \prgm_register/n837 ) );
  nand2 \prgm_register/C4337  ( .a(\prgm_register/en_not ), .b(a[418]), .out(
        \prgm_register/n838 ) );
  nand2 \prgm_register/C4338  ( .a(\prgm_register/n837 ), .b(
        \prgm_register/n838 ), .out(\prgm_register/or_signal [418]) );
  nand2 \prgm_register/C4339  ( .a(enable), .b(a[418]), .out(
        \prgm_register/n839 ) );
  nand2 \prgm_register/C4340  ( .a(\prgm_register/en_not ), .b(a[419]), .out(
        \prgm_register/n840 ) );
  nand2 \prgm_register/C4341  ( .a(\prgm_register/n839 ), .b(
        \prgm_register/n840 ), .out(\prgm_register/or_signal [419]) );
  nand2 \prgm_register/C4342  ( .a(enable), .b(a[419]), .out(
        \prgm_register/n841 ) );
  nand2 \prgm_register/C4343  ( .a(\prgm_register/en_not ), .b(a[420]), .out(
        \prgm_register/n842 ) );
  nand2 \prgm_register/C4344  ( .a(\prgm_register/n841 ), .b(
        \prgm_register/n842 ), .out(\prgm_register/or_signal [420]) );
  nand2 \prgm_register/C4345  ( .a(enable), .b(a[420]), .out(
        \prgm_register/n843 ) );
  nand2 \prgm_register/C4346  ( .a(\prgm_register/en_not ), .b(a[421]), .out(
        \prgm_register/n844 ) );
  nand2 \prgm_register/C4347  ( .a(\prgm_register/n843 ), .b(
        \prgm_register/n844 ), .out(\prgm_register/or_signal [421]) );
  nand2 \prgm_register/C4348  ( .a(enable), .b(a[421]), .out(
        \prgm_register/n845 ) );
  nand2 \prgm_register/C4349  ( .a(\prgm_register/en_not ), .b(a[422]), .out(
        \prgm_register/n846 ) );
  nand2 \prgm_register/C4350  ( .a(\prgm_register/n845 ), .b(
        \prgm_register/n846 ), .out(\prgm_register/or_signal [422]) );
  nand2 \prgm_register/C4351  ( .a(enable), .b(a[422]), .out(
        \prgm_register/n847 ) );
  nand2 \prgm_register/C4352  ( .a(\prgm_register/en_not ), .b(a[423]), .out(
        \prgm_register/n848 ) );
  nand2 \prgm_register/C4353  ( .a(\prgm_register/n847 ), .b(
        \prgm_register/n848 ), .out(\prgm_register/or_signal [423]) );
  nand2 \prgm_register/C4354  ( .a(enable), .b(a[423]), .out(
        \prgm_register/n849 ) );
  nand2 \prgm_register/C4355  ( .a(\prgm_register/en_not ), .b(a[424]), .out(
        \prgm_register/n850 ) );
  nand2 \prgm_register/C4356  ( .a(\prgm_register/n849 ), .b(
        \prgm_register/n850 ), .out(\prgm_register/or_signal [424]) );
  nand2 \prgm_register/C4357  ( .a(enable), .b(a[424]), .out(
        \prgm_register/n851 ) );
  nand2 \prgm_register/C4358  ( .a(\prgm_register/en_not ), .b(a[425]), .out(
        \prgm_register/n852 ) );
  nand2 \prgm_register/C4359  ( .a(\prgm_register/n851 ), .b(
        \prgm_register/n852 ), .out(\prgm_register/or_signal [425]) );
  nand2 \prgm_register/C4360  ( .a(enable), .b(a[425]), .out(
        \prgm_register/n853 ) );
  nand2 \prgm_register/C4361  ( .a(\prgm_register/en_not ), .b(a[426]), .out(
        \prgm_register/n854 ) );
  nand2 \prgm_register/C4362  ( .a(\prgm_register/n853 ), .b(
        \prgm_register/n854 ), .out(\prgm_register/or_signal [426]) );
  nand2 \prgm_register/C4363  ( .a(enable), .b(a[426]), .out(
        \prgm_register/n855 ) );
  nand2 \prgm_register/C4364  ( .a(\prgm_register/en_not ), .b(a[427]), .out(
        \prgm_register/n856 ) );
  nand2 \prgm_register/C4365  ( .a(\prgm_register/n855 ), .b(
        \prgm_register/n856 ), .out(\prgm_register/or_signal [427]) );
  nand2 \prgm_register/C4366  ( .a(enable), .b(a[427]), .out(
        \prgm_register/n857 ) );
  nand2 \prgm_register/C4367  ( .a(\prgm_register/en_not ), .b(a[428]), .out(
        \prgm_register/n858 ) );
  nand2 \prgm_register/C4368  ( .a(\prgm_register/n857 ), .b(
        \prgm_register/n858 ), .out(\prgm_register/or_signal [428]) );
  nand2 \prgm_register/C4369  ( .a(enable), .b(a[428]), .out(
        \prgm_register/n859 ) );
  nand2 \prgm_register/C4370  ( .a(\prgm_register/en_not ), .b(a[429]), .out(
        \prgm_register/n860 ) );
  nand2 \prgm_register/C4371  ( .a(\prgm_register/n859 ), .b(
        \prgm_register/n860 ), .out(\prgm_register/or_signal [429]) );
  nand2 \prgm_register/C4372  ( .a(enable), .b(a[429]), .out(
        \prgm_register/n861 ) );
  nand2 \prgm_register/C4373  ( .a(\prgm_register/en_not ), .b(a[430]), .out(
        \prgm_register/n862 ) );
  nand2 \prgm_register/C4374  ( .a(\prgm_register/n861 ), .b(
        \prgm_register/n862 ), .out(\prgm_register/or_signal [430]) );
  nand2 \prgm_register/C4375  ( .a(enable), .b(a[430]), .out(
        \prgm_register/n863 ) );
  nand2 \prgm_register/C4376  ( .a(\prgm_register/en_not ), .b(a[431]), .out(
        \prgm_register/n864 ) );
  nand2 \prgm_register/C4377  ( .a(\prgm_register/n863 ), .b(
        \prgm_register/n864 ), .out(\prgm_register/or_signal [431]) );
  nand2 \prgm_register/C4378  ( .a(enable), .b(a[431]), .out(
        \prgm_register/n865 ) );
  nand2 \prgm_register/C4379  ( .a(\prgm_register/en_not ), .b(a[432]), .out(
        \prgm_register/n866 ) );
  nand2 \prgm_register/C4380  ( .a(\prgm_register/n865 ), .b(
        \prgm_register/n866 ), .out(\prgm_register/or_signal [432]) );
  nand2 \prgm_register/C4381  ( .a(enable), .b(a[432]), .out(
        \prgm_register/n867 ) );
  nand2 \prgm_register/C4382  ( .a(\prgm_register/en_not ), .b(a[433]), .out(
        \prgm_register/n868 ) );
  nand2 \prgm_register/C4383  ( .a(\prgm_register/n867 ), .b(
        \prgm_register/n868 ), .out(\prgm_register/or_signal [433]) );
  nand2 \prgm_register/C4384  ( .a(enable), .b(a[433]), .out(
        \prgm_register/n869 ) );
  nand2 \prgm_register/C4385  ( .a(\prgm_register/en_not ), .b(a[434]), .out(
        \prgm_register/n870 ) );
  nand2 \prgm_register/C4386  ( .a(\prgm_register/n869 ), .b(
        \prgm_register/n870 ), .out(\prgm_register/or_signal [434]) );
  nand2 \prgm_register/C4387  ( .a(enable), .b(a[434]), .out(
        \prgm_register/n871 ) );
  nand2 \prgm_register/C4388  ( .a(\prgm_register/en_not ), .b(a[435]), .out(
        \prgm_register/n872 ) );
  nand2 \prgm_register/C4389  ( .a(\prgm_register/n871 ), .b(
        \prgm_register/n872 ), .out(\prgm_register/or_signal [435]) );
  nand2 \prgm_register/C4390  ( .a(enable), .b(a[435]), .out(
        \prgm_register/n873 ) );
  nand2 \prgm_register/C4391  ( .a(\prgm_register/en_not ), .b(a[436]), .out(
        \prgm_register/n874 ) );
  nand2 \prgm_register/C4392  ( .a(\prgm_register/n873 ), .b(
        \prgm_register/n874 ), .out(\prgm_register/or_signal [436]) );
  nand2 \prgm_register/C4393  ( .a(enable), .b(a[436]), .out(
        \prgm_register/n875 ) );
  nand2 \prgm_register/C4394  ( .a(\prgm_register/en_not ), .b(a[437]), .out(
        \prgm_register/n876 ) );
  nand2 \prgm_register/C4395  ( .a(\prgm_register/n875 ), .b(
        \prgm_register/n876 ), .out(\prgm_register/or_signal [437]) );
  nand2 \prgm_register/C4396  ( .a(enable), .b(a[437]), .out(
        \prgm_register/n877 ) );
  nand2 \prgm_register/C4397  ( .a(\prgm_register/en_not ), .b(a[438]), .out(
        \prgm_register/n878 ) );
  nand2 \prgm_register/C4398  ( .a(\prgm_register/n877 ), .b(
        \prgm_register/n878 ), .out(\prgm_register/or_signal [438]) );
  nand2 \prgm_register/C4399  ( .a(enable), .b(a[438]), .out(
        \prgm_register/n879 ) );
  nand2 \prgm_register/C4400  ( .a(\prgm_register/en_not ), .b(a[439]), .out(
        \prgm_register/n880 ) );
  nand2 \prgm_register/C4401  ( .a(\prgm_register/n879 ), .b(
        \prgm_register/n880 ), .out(\prgm_register/or_signal [439]) );
  nand2 \prgm_register/C4402  ( .a(enable), .b(a[439]), .out(
        \prgm_register/n881 ) );
  nand2 \prgm_register/C4403  ( .a(\prgm_register/en_not ), .b(a[440]), .out(
        \prgm_register/n882 ) );
  nand2 \prgm_register/C4404  ( .a(\prgm_register/n881 ), .b(
        \prgm_register/n882 ), .out(\prgm_register/or_signal [440]) );
  nand2 \prgm_register/C4405  ( .a(enable), .b(a[440]), .out(
        \prgm_register/n883 ) );
  nand2 \prgm_register/C4406  ( .a(\prgm_register/en_not ), .b(a[441]), .out(
        \prgm_register/n884 ) );
  nand2 \prgm_register/C4407  ( .a(\prgm_register/n883 ), .b(
        \prgm_register/n884 ), .out(\prgm_register/or_signal [441]) );
  nand2 \prgm_register/C4408  ( .a(enable), .b(a[441]), .out(
        \prgm_register/n885 ) );
  nand2 \prgm_register/C4409  ( .a(\prgm_register/en_not ), .b(a[442]), .out(
        \prgm_register/n886 ) );
  nand2 \prgm_register/C4410  ( .a(\prgm_register/n885 ), .b(
        \prgm_register/n886 ), .out(\prgm_register/or_signal [442]) );
  nand2 \prgm_register/C4411  ( .a(enable), .b(a[442]), .out(
        \prgm_register/n887 ) );
  nand2 \prgm_register/C4412  ( .a(\prgm_register/en_not ), .b(a[443]), .out(
        \prgm_register/n888 ) );
  nand2 \prgm_register/C4413  ( .a(\prgm_register/n887 ), .b(
        \prgm_register/n888 ), .out(\prgm_register/or_signal [443]) );
  nand2 \prgm_register/C4414  ( .a(enable), .b(a[443]), .out(
        \prgm_register/n889 ) );
  nand2 \prgm_register/C4415  ( .a(\prgm_register/en_not ), .b(a[444]), .out(
        \prgm_register/n890 ) );
  nand2 \prgm_register/C4416  ( .a(\prgm_register/n889 ), .b(
        \prgm_register/n890 ), .out(\prgm_register/or_signal [444]) );
  nand2 \prgm_register/C4417  ( .a(enable), .b(a[444]), .out(
        \prgm_register/n891 ) );
  nand2 \prgm_register/C4418  ( .a(\prgm_register/en_not ), .b(a[445]), .out(
        \prgm_register/n892 ) );
  nand2 \prgm_register/C4419  ( .a(\prgm_register/n891 ), .b(
        \prgm_register/n892 ), .out(\prgm_register/or_signal [445]) );
  nand2 \prgm_register/C4420  ( .a(enable), .b(a[445]), .out(
        \prgm_register/n893 ) );
  nand2 \prgm_register/C4421  ( .a(\prgm_register/en_not ), .b(a[446]), .out(
        \prgm_register/n894 ) );
  nand2 \prgm_register/C4422  ( .a(\prgm_register/n893 ), .b(
        \prgm_register/n894 ), .out(\prgm_register/or_signal [446]) );
  nand2 \prgm_register/C4423  ( .a(enable), .b(a[446]), .out(
        \prgm_register/n895 ) );
  nand2 \prgm_register/C4424  ( .a(\prgm_register/en_not ), .b(a[447]), .out(
        \prgm_register/n896 ) );
  nand2 \prgm_register/C4425  ( .a(\prgm_register/n895 ), .b(
        \prgm_register/n896 ), .out(\prgm_register/or_signal [447]) );
  nand2 \prgm_register/C4426  ( .a(enable), .b(a[447]), .out(
        \prgm_register/n897 ) );
  nand2 \prgm_register/C4427  ( .a(\prgm_register/en_not ), .b(a[448]), .out(
        \prgm_register/n898 ) );
  nand2 \prgm_register/C4428  ( .a(\prgm_register/n897 ), .b(
        \prgm_register/n898 ), .out(\prgm_register/or_signal [448]) );
  nand2 \prgm_register/C4429  ( .a(enable), .b(a[448]), .out(
        \prgm_register/n899 ) );
  nand2 \prgm_register/C4430  ( .a(\prgm_register/en_not ), .b(a[449]), .out(
        \prgm_register/n900 ) );
  nand2 \prgm_register/C4431  ( .a(\prgm_register/n899 ), .b(
        \prgm_register/n900 ), .out(\prgm_register/or_signal [449]) );
  nand2 \prgm_register/C4432  ( .a(enable), .b(a[449]), .out(
        \prgm_register/n901 ) );
  nand2 \prgm_register/C4433  ( .a(\prgm_register/en_not ), .b(a[450]), .out(
        \prgm_register/n902 ) );
  nand2 \prgm_register/C4434  ( .a(\prgm_register/n901 ), .b(
        \prgm_register/n902 ), .out(\prgm_register/or_signal [450]) );
  nand2 \prgm_register/C4435  ( .a(enable), .b(a[450]), .out(
        \prgm_register/n903 ) );
  nand2 \prgm_register/C4436  ( .a(\prgm_register/en_not ), .b(a[451]), .out(
        \prgm_register/n904 ) );
  nand2 \prgm_register/C4437  ( .a(\prgm_register/n903 ), .b(
        \prgm_register/n904 ), .out(\prgm_register/or_signal [451]) );
  nand2 \prgm_register/C4438  ( .a(enable), .b(a[451]), .out(
        \prgm_register/n905 ) );
  nand2 \prgm_register/C4439  ( .a(\prgm_register/en_not ), .b(a[452]), .out(
        \prgm_register/n906 ) );
  nand2 \prgm_register/C4440  ( .a(\prgm_register/n905 ), .b(
        \prgm_register/n906 ), .out(\prgm_register/or_signal [452]) );
  nand2 \prgm_register/C4441  ( .a(enable), .b(a[452]), .out(
        \prgm_register/n907 ) );
  nand2 \prgm_register/C4442  ( .a(\prgm_register/en_not ), .b(a[453]), .out(
        \prgm_register/n908 ) );
  nand2 \prgm_register/C4443  ( .a(\prgm_register/n907 ), .b(
        \prgm_register/n908 ), .out(\prgm_register/or_signal [453]) );
  nand2 \prgm_register/C4444  ( .a(enable), .b(a[453]), .out(
        \prgm_register/n909 ) );
  nand2 \prgm_register/C4445  ( .a(\prgm_register/en_not ), .b(a[454]), .out(
        \prgm_register/n910 ) );
  nand2 \prgm_register/C4446  ( .a(\prgm_register/n909 ), .b(
        \prgm_register/n910 ), .out(\prgm_register/or_signal [454]) );
  nand2 \prgm_register/C4447  ( .a(enable), .b(a[454]), .out(
        \prgm_register/n911 ) );
  nand2 \prgm_register/C4448  ( .a(\prgm_register/en_not ), .b(a[455]), .out(
        \prgm_register/n912 ) );
  nand2 \prgm_register/C4449  ( .a(\prgm_register/n911 ), .b(
        \prgm_register/n912 ), .out(\prgm_register/or_signal [455]) );
  nand2 \prgm_register/C4450  ( .a(enable), .b(a[455]), .out(
        \prgm_register/n913 ) );
  nand2 \prgm_register/C4451  ( .a(\prgm_register/en_not ), .b(a[456]), .out(
        \prgm_register/n914 ) );
  nand2 \prgm_register/C4452  ( .a(\prgm_register/n913 ), .b(
        \prgm_register/n914 ), .out(\prgm_register/or_signal [456]) );
  nand2 \prgm_register/C4453  ( .a(enable), .b(a[456]), .out(
        \prgm_register/n915 ) );
  nand2 \prgm_register/C4454  ( .a(\prgm_register/en_not ), .b(a[457]), .out(
        \prgm_register/n916 ) );
  nand2 \prgm_register/C4455  ( .a(\prgm_register/n915 ), .b(
        \prgm_register/n916 ), .out(\prgm_register/or_signal [457]) );
  nand2 \prgm_register/C4456  ( .a(enable), .b(a[457]), .out(
        \prgm_register/n917 ) );
  nand2 \prgm_register/C4457  ( .a(\prgm_register/en_not ), .b(a[458]), .out(
        \prgm_register/n918 ) );
  nand2 \prgm_register/C4458  ( .a(\prgm_register/n917 ), .b(
        \prgm_register/n918 ), .out(\prgm_register/or_signal [458]) );
  nand2 \prgm_register/C4459  ( .a(enable), .b(a[458]), .out(
        \prgm_register/n919 ) );
  nand2 \prgm_register/C4460  ( .a(\prgm_register/en_not ), .b(a[459]), .out(
        \prgm_register/n920 ) );
  nand2 \prgm_register/C4461  ( .a(\prgm_register/n919 ), .b(
        \prgm_register/n920 ), .out(\prgm_register/or_signal [459]) );
  nand2 \prgm_register/C4462  ( .a(enable), .b(a[459]), .out(
        \prgm_register/n921 ) );
  nand2 \prgm_register/C4463  ( .a(\prgm_register/en_not ), .b(a[460]), .out(
        \prgm_register/n922 ) );
  nand2 \prgm_register/C4464  ( .a(\prgm_register/n921 ), .b(
        \prgm_register/n922 ), .out(\prgm_register/or_signal [460]) );
  nand2 \prgm_register/C4465  ( .a(enable), .b(a[460]), .out(
        \prgm_register/n923 ) );
  nand2 \prgm_register/C4466  ( .a(\prgm_register/en_not ), .b(a[461]), .out(
        \prgm_register/n924 ) );
  nand2 \prgm_register/C4467  ( .a(\prgm_register/n923 ), .b(
        \prgm_register/n924 ), .out(\prgm_register/or_signal [461]) );
  nand2 \prgm_register/C4468  ( .a(enable), .b(a[461]), .out(
        \prgm_register/n925 ) );
  nand2 \prgm_register/C4469  ( .a(\prgm_register/en_not ), .b(a[462]), .out(
        \prgm_register/n926 ) );
  nand2 \prgm_register/C4470  ( .a(\prgm_register/n925 ), .b(
        \prgm_register/n926 ), .out(\prgm_register/or_signal [462]) );
  nand2 \prgm_register/C4471  ( .a(enable), .b(a[462]), .out(
        \prgm_register/n927 ) );
  nand2 \prgm_register/C4472  ( .a(\prgm_register/en_not ), .b(a[463]), .out(
        \prgm_register/n928 ) );
  nand2 \prgm_register/C4473  ( .a(\prgm_register/n927 ), .b(
        \prgm_register/n928 ), .out(\prgm_register/or_signal [463]) );
  nand2 \prgm_register/C4474  ( .a(enable), .b(a[463]), .out(
        \prgm_register/n929 ) );
  nand2 \prgm_register/C4475  ( .a(\prgm_register/en_not ), .b(a[464]), .out(
        \prgm_register/n930 ) );
  nand2 \prgm_register/C4476  ( .a(\prgm_register/n929 ), .b(
        \prgm_register/n930 ), .out(\prgm_register/or_signal [464]) );
  nand2 \prgm_register/C4477  ( .a(enable), .b(a[464]), .out(
        \prgm_register/n931 ) );
  nand2 \prgm_register/C4478  ( .a(\prgm_register/en_not ), .b(a[465]), .out(
        \prgm_register/n932 ) );
  nand2 \prgm_register/C4479  ( .a(\prgm_register/n931 ), .b(
        \prgm_register/n932 ), .out(\prgm_register/or_signal [465]) );
  nand2 \prgm_register/C4480  ( .a(enable), .b(a[465]), .out(
        \prgm_register/n933 ) );
  nand2 \prgm_register/C4481  ( .a(\prgm_register/en_not ), .b(a[466]), .out(
        \prgm_register/n934 ) );
  nand2 \prgm_register/C4482  ( .a(\prgm_register/n933 ), .b(
        \prgm_register/n934 ), .out(\prgm_register/or_signal [466]) );
  nand2 \prgm_register/C4483  ( .a(enable), .b(a[466]), .out(
        \prgm_register/n935 ) );
  nand2 \prgm_register/C4484  ( .a(\prgm_register/en_not ), .b(a[467]), .out(
        \prgm_register/n936 ) );
  nand2 \prgm_register/C4485  ( .a(\prgm_register/n935 ), .b(
        \prgm_register/n936 ), .out(\prgm_register/or_signal [467]) );
  nand2 \prgm_register/C4486  ( .a(enable), .b(a[467]), .out(
        \prgm_register/n937 ) );
  nand2 \prgm_register/C4487  ( .a(\prgm_register/en_not ), .b(a[468]), .out(
        \prgm_register/n938 ) );
  nand2 \prgm_register/C4488  ( .a(\prgm_register/n937 ), .b(
        \prgm_register/n938 ), .out(\prgm_register/or_signal [468]) );
  nand2 \prgm_register/C4489  ( .a(enable), .b(a[468]), .out(
        \prgm_register/n939 ) );
  nand2 \prgm_register/C4490  ( .a(\prgm_register/en_not ), .b(a[469]), .out(
        \prgm_register/n940 ) );
  nand2 \prgm_register/C4491  ( .a(\prgm_register/n939 ), .b(
        \prgm_register/n940 ), .out(\prgm_register/or_signal [469]) );
  nand2 \prgm_register/C4492  ( .a(enable), .b(a[469]), .out(
        \prgm_register/n941 ) );
  nand2 \prgm_register/C4493  ( .a(\prgm_register/en_not ), .b(a[470]), .out(
        \prgm_register/n942 ) );
  nand2 \prgm_register/C4494  ( .a(\prgm_register/n941 ), .b(
        \prgm_register/n942 ), .out(\prgm_register/or_signal [470]) );
  nand2 \prgm_register/C4495  ( .a(enable), .b(a[470]), .out(
        \prgm_register/n943 ) );
  nand2 \prgm_register/C4496  ( .a(\prgm_register/en_not ), .b(a[471]), .out(
        \prgm_register/n944 ) );
  nand2 \prgm_register/C4497  ( .a(\prgm_register/n943 ), .b(
        \prgm_register/n944 ), .out(\prgm_register/or_signal [471]) );
  nand2 \prgm_register/C4498  ( .a(enable), .b(a[471]), .out(
        \prgm_register/n945 ) );
  nand2 \prgm_register/C4499  ( .a(\prgm_register/en_not ), .b(a[472]), .out(
        \prgm_register/n946 ) );
  nand2 \prgm_register/C4500  ( .a(\prgm_register/n945 ), .b(
        \prgm_register/n946 ), .out(\prgm_register/or_signal [472]) );
  nand2 \prgm_register/C4501  ( .a(enable), .b(a[472]), .out(
        \prgm_register/n947 ) );
  nand2 \prgm_register/C4502  ( .a(\prgm_register/en_not ), .b(a[473]), .out(
        \prgm_register/n948 ) );
  nand2 \prgm_register/C4503  ( .a(\prgm_register/n947 ), .b(
        \prgm_register/n948 ), .out(\prgm_register/or_signal [473]) );
  nand2 \prgm_register/C4504  ( .a(enable), .b(a[473]), .out(
        \prgm_register/n949 ) );
  nand2 \prgm_register/C4505  ( .a(\prgm_register/en_not ), .b(a[474]), .out(
        \prgm_register/n950 ) );
  nand2 \prgm_register/C4506  ( .a(\prgm_register/n949 ), .b(
        \prgm_register/n950 ), .out(\prgm_register/or_signal [474]) );
  nand2 \prgm_register/C4507  ( .a(enable), .b(a[474]), .out(
        \prgm_register/n951 ) );
  nand2 \prgm_register/C4508  ( .a(\prgm_register/en_not ), .b(a[475]), .out(
        \prgm_register/n952 ) );
  nand2 \prgm_register/C4509  ( .a(\prgm_register/n951 ), .b(
        \prgm_register/n952 ), .out(\prgm_register/or_signal [475]) );
  nand2 \prgm_register/C4510  ( .a(enable), .b(a[475]), .out(
        \prgm_register/n953 ) );
  nand2 \prgm_register/C4511  ( .a(\prgm_register/en_not ), .b(a[476]), .out(
        \prgm_register/n954 ) );
  nand2 \prgm_register/C4512  ( .a(\prgm_register/n953 ), .b(
        \prgm_register/n954 ), .out(\prgm_register/or_signal [476]) );
  nand2 \prgm_register/C4513  ( .a(enable), .b(a[476]), .out(
        \prgm_register/n955 ) );
  nand2 \prgm_register/C4514  ( .a(\prgm_register/en_not ), .b(a[477]), .out(
        \prgm_register/n956 ) );
  nand2 \prgm_register/C4515  ( .a(\prgm_register/n955 ), .b(
        \prgm_register/n956 ), .out(\prgm_register/or_signal [477]) );
  nand2 \prgm_register/C4516  ( .a(enable), .b(a[477]), .out(
        \prgm_register/n957 ) );
  nand2 \prgm_register/C4517  ( .a(\prgm_register/en_not ), .b(a[478]), .out(
        \prgm_register/n958 ) );
  nand2 \prgm_register/C4518  ( .a(\prgm_register/n957 ), .b(
        \prgm_register/n958 ), .out(\prgm_register/or_signal [478]) );
  nand2 \prgm_register/C4519  ( .a(enable), .b(a[478]), .out(
        \prgm_register/n959 ) );
  nand2 \prgm_register/C4520  ( .a(\prgm_register/en_not ), .b(a[479]), .out(
        \prgm_register/n960 ) );
  nand2 \prgm_register/C4521  ( .a(\prgm_register/n959 ), .b(
        \prgm_register/n960 ), .out(\prgm_register/or_signal [479]) );
  nand2 \prgm_register/C4522  ( .a(enable), .b(a[479]), .out(
        \prgm_register/n961 ) );
  nand2 \prgm_register/C4523  ( .a(\prgm_register/en_not ), .b(a[480]), .out(
        \prgm_register/n962 ) );
  nand2 \prgm_register/C4524  ( .a(\prgm_register/n961 ), .b(
        \prgm_register/n962 ), .out(\prgm_register/or_signal [480]) );
  nand2 \prgm_register/C4525  ( .a(enable), .b(a[480]), .out(
        \prgm_register/n963 ) );
  nand2 \prgm_register/C4526  ( .a(\prgm_register/en_not ), .b(a[481]), .out(
        \prgm_register/n964 ) );
  nand2 \prgm_register/C4527  ( .a(\prgm_register/n963 ), .b(
        \prgm_register/n964 ), .out(\prgm_register/or_signal [481]) );
  nand2 \prgm_register/C4528  ( .a(enable), .b(a[481]), .out(
        \prgm_register/n965 ) );
  nand2 \prgm_register/C4529  ( .a(\prgm_register/en_not ), .b(a[482]), .out(
        \prgm_register/n966 ) );
  nand2 \prgm_register/C4530  ( .a(\prgm_register/n965 ), .b(
        \prgm_register/n966 ), .out(\prgm_register/or_signal [482]) );
  nand2 \prgm_register/C4531  ( .a(enable), .b(a[482]), .out(
        \prgm_register/n967 ) );
  nand2 \prgm_register/C4532  ( .a(\prgm_register/en_not ), .b(a[483]), .out(
        \prgm_register/n968 ) );
  nand2 \prgm_register/C4533  ( .a(\prgm_register/n967 ), .b(
        \prgm_register/n968 ), .out(\prgm_register/or_signal [483]) );
  nand2 \prgm_register/C4534  ( .a(enable), .b(a[483]), .out(
        \prgm_register/n969 ) );
  nand2 \prgm_register/C4535  ( .a(\prgm_register/en_not ), .b(a[484]), .out(
        \prgm_register/n970 ) );
  nand2 \prgm_register/C4536  ( .a(\prgm_register/n969 ), .b(
        \prgm_register/n970 ), .out(\prgm_register/or_signal [484]) );
  nand2 \prgm_register/C4537  ( .a(enable), .b(a[484]), .out(
        \prgm_register/n971 ) );
  nand2 \prgm_register/C4538  ( .a(\prgm_register/en_not ), .b(a[485]), .out(
        \prgm_register/n972 ) );
  nand2 \prgm_register/C4539  ( .a(\prgm_register/n971 ), .b(
        \prgm_register/n972 ), .out(\prgm_register/or_signal [485]) );
  nand2 \prgm_register/C4540  ( .a(enable), .b(a[485]), .out(
        \prgm_register/n973 ) );
  nand2 \prgm_register/C4541  ( .a(\prgm_register/en_not ), .b(a[486]), .out(
        \prgm_register/n974 ) );
  nand2 \prgm_register/C4542  ( .a(\prgm_register/n973 ), .b(
        \prgm_register/n974 ), .out(\prgm_register/or_signal [486]) );
  nand2 \prgm_register/C4543  ( .a(enable), .b(a[486]), .out(
        \prgm_register/n975 ) );
  nand2 \prgm_register/C4544  ( .a(\prgm_register/en_not ), .b(a[487]), .out(
        \prgm_register/n976 ) );
  nand2 \prgm_register/C4545  ( .a(\prgm_register/n975 ), .b(
        \prgm_register/n976 ), .out(\prgm_register/or_signal [487]) );
  nand2 \prgm_register/C4546  ( .a(enable), .b(a[487]), .out(
        \prgm_register/n977 ) );
  nand2 \prgm_register/C4547  ( .a(\prgm_register/en_not ), .b(a[488]), .out(
        \prgm_register/n978 ) );
  nand2 \prgm_register/C4548  ( .a(\prgm_register/n977 ), .b(
        \prgm_register/n978 ), .out(\prgm_register/or_signal [488]) );
  nand2 \prgm_register/C4549  ( .a(enable), .b(a[488]), .out(
        \prgm_register/n979 ) );
  nand2 \prgm_register/C4550  ( .a(\prgm_register/en_not ), .b(a[489]), .out(
        \prgm_register/n980 ) );
  nand2 \prgm_register/C4551  ( .a(\prgm_register/n979 ), .b(
        \prgm_register/n980 ), .out(\prgm_register/or_signal [489]) );
  nand2 \prgm_register/C4552  ( .a(enable), .b(a[489]), .out(
        \prgm_register/n981 ) );
  nand2 \prgm_register/C4553  ( .a(\prgm_register/en_not ), .b(a[490]), .out(
        \prgm_register/n982 ) );
  nand2 \prgm_register/C4554  ( .a(\prgm_register/n981 ), .b(
        \prgm_register/n982 ), .out(\prgm_register/or_signal [490]) );
  nand2 \prgm_register/C4555  ( .a(enable), .b(a[490]), .out(
        \prgm_register/n983 ) );
  nand2 \prgm_register/C4556  ( .a(\prgm_register/en_not ), .b(a[491]), .out(
        \prgm_register/n984 ) );
  nand2 \prgm_register/C4557  ( .a(\prgm_register/n983 ), .b(
        \prgm_register/n984 ), .out(\prgm_register/or_signal [491]) );
  nand2 \prgm_register/C4558  ( .a(enable), .b(a[491]), .out(
        \prgm_register/n985 ) );
  nand2 \prgm_register/C4559  ( .a(\prgm_register/en_not ), .b(a[492]), .out(
        \prgm_register/n986 ) );
  nand2 \prgm_register/C4560  ( .a(\prgm_register/n985 ), .b(
        \prgm_register/n986 ), .out(\prgm_register/or_signal [492]) );
  nand2 \prgm_register/C4561  ( .a(enable), .b(a[492]), .out(
        \prgm_register/n987 ) );
  nand2 \prgm_register/C4562  ( .a(\prgm_register/en_not ), .b(a[493]), .out(
        \prgm_register/n988 ) );
  nand2 \prgm_register/C4563  ( .a(\prgm_register/n987 ), .b(
        \prgm_register/n988 ), .out(\prgm_register/or_signal [493]) );
  nand2 \prgm_register/C4564  ( .a(enable), .b(a[493]), .out(
        \prgm_register/n989 ) );
  nand2 \prgm_register/C4565  ( .a(\prgm_register/en_not ), .b(a[494]), .out(
        \prgm_register/n990 ) );
  nand2 \prgm_register/C4566  ( .a(\prgm_register/n989 ), .b(
        \prgm_register/n990 ), .out(\prgm_register/or_signal [494]) );
  nand2 \prgm_register/C4567  ( .a(enable), .b(a[494]), .out(
        \prgm_register/n991 ) );
  nand2 \prgm_register/C4568  ( .a(\prgm_register/en_not ), .b(a[495]), .out(
        \prgm_register/n992 ) );
  nand2 \prgm_register/C4569  ( .a(\prgm_register/n991 ), .b(
        \prgm_register/n992 ), .out(\prgm_register/or_signal [495]) );
  nand2 \prgm_register/C4570  ( .a(enable), .b(a[495]), .out(
        \prgm_register/n993 ) );
  nand2 \prgm_register/C4571  ( .a(\prgm_register/en_not ), .b(a[496]), .out(
        \prgm_register/n994 ) );
  nand2 \prgm_register/C4572  ( .a(\prgm_register/n993 ), .b(
        \prgm_register/n994 ), .out(\prgm_register/or_signal [496]) );
  nand2 \prgm_register/C4573  ( .a(enable), .b(a[496]), .out(
        \prgm_register/n995 ) );
  nand2 \prgm_register/C4574  ( .a(\prgm_register/en_not ), .b(a[497]), .out(
        \prgm_register/n996 ) );
  nand2 \prgm_register/C4575  ( .a(\prgm_register/n995 ), .b(
        \prgm_register/n996 ), .out(\prgm_register/or_signal [497]) );
  nand2 \prgm_register/C4576  ( .a(enable), .b(a[497]), .out(
        \prgm_register/n997 ) );
  nand2 \prgm_register/C4577  ( .a(\prgm_register/en_not ), .b(a[498]), .out(
        \prgm_register/n998 ) );
  nand2 \prgm_register/C4578  ( .a(\prgm_register/n997 ), .b(
        \prgm_register/n998 ), .out(\prgm_register/or_signal [498]) );
  nand2 \prgm_register/C4579  ( .a(enable), .b(a[498]), .out(
        \prgm_register/n999 ) );
  nand2 \prgm_register/C4580  ( .a(\prgm_register/en_not ), .b(a[499]), .out(
        \prgm_register/n1000 ) );
  nand2 \prgm_register/C4581  ( .a(\prgm_register/n999 ), .b(
        \prgm_register/n1000 ), .out(\prgm_register/or_signal [499]) );
  nand2 \prgm_register/C4582  ( .a(enable), .b(a[499]), .out(
        \prgm_register/n1001 ) );
  nand2 \prgm_register/C4583  ( .a(\prgm_register/en_not ), .b(a[500]), .out(
        \prgm_register/n1002 ) );
  nand2 \prgm_register/C4584  ( .a(\prgm_register/n1001 ), .b(
        \prgm_register/n1002 ), .out(\prgm_register/or_signal [500]) );
  nand2 \prgm_register/C4585  ( .a(enable), .b(a[500]), .out(
        \prgm_register/n1003 ) );
  nand2 \prgm_register/C4586  ( .a(\prgm_register/en_not ), .b(a[501]), .out(
        \prgm_register/n1004 ) );
  nand2 \prgm_register/C4587  ( .a(\prgm_register/n1003 ), .b(
        \prgm_register/n1004 ), .out(\prgm_register/or_signal [501]) );
  nand2 \prgm_register/C4588  ( .a(enable), .b(a[501]), .out(
        \prgm_register/n1005 ) );
  nand2 \prgm_register/C4589  ( .a(\prgm_register/en_not ), .b(a[502]), .out(
        \prgm_register/n1006 ) );
  nand2 \prgm_register/C4590  ( .a(\prgm_register/n1005 ), .b(
        \prgm_register/n1006 ), .out(\prgm_register/or_signal [502]) );
  nand2 \prgm_register/C4591  ( .a(enable), .b(a[502]), .out(
        \prgm_register/n1007 ) );
  nand2 \prgm_register/C4592  ( .a(\prgm_register/en_not ), .b(a[503]), .out(
        \prgm_register/n1008 ) );
  nand2 \prgm_register/C4593  ( .a(\prgm_register/n1007 ), .b(
        \prgm_register/n1008 ), .out(\prgm_register/or_signal [503]) );
  nand2 \prgm_register/C4594  ( .a(enable), .b(a[503]), .out(
        \prgm_register/n1009 ) );
  nand2 \prgm_register/C4595  ( .a(\prgm_register/en_not ), .b(a[504]), .out(
        \prgm_register/n1010 ) );
  nand2 \prgm_register/C4596  ( .a(\prgm_register/n1009 ), .b(
        \prgm_register/n1010 ), .out(\prgm_register/or_signal [504]) );
  nand2 \prgm_register/C4597  ( .a(enable), .b(a[504]), .out(
        \prgm_register/n1011 ) );
  nand2 \prgm_register/C4598  ( .a(\prgm_register/en_not ), .b(a[505]), .out(
        \prgm_register/n1012 ) );
  nand2 \prgm_register/C4599  ( .a(\prgm_register/n1011 ), .b(
        \prgm_register/n1012 ), .out(\prgm_register/or_signal [505]) );
  nand2 \prgm_register/C4600  ( .a(enable), .b(a[505]), .out(
        \prgm_register/n1013 ) );
  nand2 \prgm_register/C4601  ( .a(\prgm_register/en_not ), .b(a[506]), .out(
        \prgm_register/n1014 ) );
  nand2 \prgm_register/C4602  ( .a(\prgm_register/n1013 ), .b(
        \prgm_register/n1014 ), .out(\prgm_register/or_signal [506]) );
  nand2 \prgm_register/C4603  ( .a(enable), .b(a[506]), .out(
        \prgm_register/n1015 ) );
  nand2 \prgm_register/C4604  ( .a(\prgm_register/en_not ), .b(a[507]), .out(
        \prgm_register/n1016 ) );
  nand2 \prgm_register/C4605  ( .a(\prgm_register/n1015 ), .b(
        \prgm_register/n1016 ), .out(\prgm_register/or_signal [507]) );
  nand2 \prgm_register/C4606  ( .a(enable), .b(a[507]), .out(
        \prgm_register/n1017 ) );
  nand2 \prgm_register/C4607  ( .a(\prgm_register/en_not ), .b(a[508]), .out(
        \prgm_register/n1018 ) );
  nand2 \prgm_register/C4608  ( .a(\prgm_register/n1017 ), .b(
        \prgm_register/n1018 ), .out(\prgm_register/or_signal [508]) );
  nand2 \prgm_register/C4609  ( .a(enable), .b(a[508]), .out(
        \prgm_register/n1019 ) );
  nand2 \prgm_register/C4610  ( .a(\prgm_register/en_not ), .b(a[509]), .out(
        \prgm_register/n1020 ) );
  nand2 \prgm_register/C4611  ( .a(\prgm_register/n1019 ), .b(
        \prgm_register/n1020 ), .out(\prgm_register/or_signal [509]) );
  nand2 \prgm_register/C4612  ( .a(enable), .b(a[509]), .out(
        \prgm_register/n1021 ) );
  nand2 \prgm_register/C4613  ( .a(\prgm_register/en_not ), .b(a[510]), .out(
        \prgm_register/n1022 ) );
  nand2 \prgm_register/C4614  ( .a(\prgm_register/n1021 ), .b(
        \prgm_register/n1022 ), .out(\prgm_register/or_signal [510]) );
  nand2 \prgm_register/C4615  ( .a(enable), .b(a[510]), .out(
        \prgm_register/n1023 ) );
  nand2 \prgm_register/C4616  ( .a(\prgm_register/en_not ), .b(a[511]), .out(
        \prgm_register/n1024 ) );
  nand2 \prgm_register/C4617  ( .a(\prgm_register/n1023 ), .b(
        \prgm_register/n1024 ), .out(\prgm_register/or_signal [511]) );
  nand2 \prgm_register/C4618  ( .a(enable), .b(a[511]), .out(
        \prgm_register/n1025 ) );
  nand2 \prgm_register/C4619  ( .a(\prgm_register/en_not ), .b(a[512]), .out(
        \prgm_register/n1026 ) );
  nand2 \prgm_register/C4620  ( .a(\prgm_register/n1025 ), .b(
        \prgm_register/n1026 ), .out(\prgm_register/or_signal [512]) );
  nand2 \prgm_register/C4621  ( .a(enable), .b(a[512]), .out(
        \prgm_register/n1027 ) );
  nand2 \prgm_register/C4622  ( .a(\prgm_register/en_not ), .b(a[513]), .out(
        \prgm_register/n1028 ) );
  nand2 \prgm_register/C4623  ( .a(\prgm_register/n1027 ), .b(
        \prgm_register/n1028 ), .out(\prgm_register/or_signal [513]) );
  nand2 \prgm_register/C4624  ( .a(enable), .b(a[513]), .out(
        \prgm_register/n1029 ) );
  nand2 \prgm_register/C4625  ( .a(\prgm_register/en_not ), .b(a[514]), .out(
        \prgm_register/n1030 ) );
  nand2 \prgm_register/C4626  ( .a(\prgm_register/n1029 ), .b(
        \prgm_register/n1030 ), .out(\prgm_register/or_signal [514]) );
  nand2 \prgm_register/C4627  ( .a(enable), .b(a[514]), .out(
        \prgm_register/n1031 ) );
  nand2 \prgm_register/C4628  ( .a(\prgm_register/en_not ), .b(a[515]), .out(
        \prgm_register/n1032 ) );
  nand2 \prgm_register/C4629  ( .a(\prgm_register/n1031 ), .b(
        \prgm_register/n1032 ), .out(\prgm_register/or_signal [515]) );
  nand2 \prgm_register/C4630  ( .a(enable), .b(a[515]), .out(
        \prgm_register/n1033 ) );
  nand2 \prgm_register/C4631  ( .a(\prgm_register/en_not ), .b(a[516]), .out(
        \prgm_register/n1034 ) );
  nand2 \prgm_register/C4632  ( .a(\prgm_register/n1033 ), .b(
        \prgm_register/n1034 ), .out(\prgm_register/or_signal [516]) );
  nand2 \prgm_register/C4633  ( .a(enable), .b(a[516]), .out(
        \prgm_register/n1035 ) );
  nand2 \prgm_register/C4634  ( .a(\prgm_register/en_not ), .b(a[517]), .out(
        \prgm_register/n1036 ) );
  nand2 \prgm_register/C4635  ( .a(\prgm_register/n1035 ), .b(
        \prgm_register/n1036 ), .out(\prgm_register/or_signal [517]) );
  nand2 \prgm_register/C4636  ( .a(enable), .b(a[517]), .out(
        \prgm_register/n1037 ) );
  nand2 \prgm_register/C4637  ( .a(\prgm_register/en_not ), .b(a[518]), .out(
        \prgm_register/n1038 ) );
  nand2 \prgm_register/C4638  ( .a(\prgm_register/n1037 ), .b(
        \prgm_register/n1038 ), .out(\prgm_register/or_signal [518]) );
  nand2 \prgm_register/C4639  ( .a(enable), .b(a[518]), .out(
        \prgm_register/n1039 ) );
  nand2 \prgm_register/C4640  ( .a(\prgm_register/en_not ), .b(a[519]), .out(
        \prgm_register/n1040 ) );
  nand2 \prgm_register/C4641  ( .a(\prgm_register/n1039 ), .b(
        \prgm_register/n1040 ), .out(\prgm_register/or_signal [519]) );
  nand2 \prgm_register/C4642  ( .a(enable), .b(a[519]), .out(
        \prgm_register/n1041 ) );
  nand2 \prgm_register/C4643  ( .a(\prgm_register/en_not ), .b(a[520]), .out(
        \prgm_register/n1042 ) );
  nand2 \prgm_register/C4644  ( .a(\prgm_register/n1041 ), .b(
        \prgm_register/n1042 ), .out(\prgm_register/or_signal [520]) );
  nand2 \prgm_register/C4645  ( .a(enable), .b(a[520]), .out(
        \prgm_register/n1043 ) );
  nand2 \prgm_register/C4646  ( .a(\prgm_register/en_not ), .b(a[521]), .out(
        \prgm_register/n1044 ) );
  nand2 \prgm_register/C4647  ( .a(\prgm_register/n1043 ), .b(
        \prgm_register/n1044 ), .out(\prgm_register/or_signal [521]) );
  nand2 \prgm_register/C4648  ( .a(enable), .b(a[521]), .out(
        \prgm_register/n1045 ) );
  nand2 \prgm_register/C4649  ( .a(\prgm_register/en_not ), .b(a[522]), .out(
        \prgm_register/n1046 ) );
  nand2 \prgm_register/C4650  ( .a(\prgm_register/n1045 ), .b(
        \prgm_register/n1046 ), .out(\prgm_register/or_signal [522]) );
  nand2 \prgm_register/C4651  ( .a(enable), .b(a[522]), .out(
        \prgm_register/n1047 ) );
  nand2 \prgm_register/C4652  ( .a(\prgm_register/en_not ), .b(a[523]), .out(
        \prgm_register/n1048 ) );
  nand2 \prgm_register/C4653  ( .a(\prgm_register/n1047 ), .b(
        \prgm_register/n1048 ), .out(\prgm_register/or_signal [523]) );
  nand2 \prgm_register/C4654  ( .a(enable), .b(a[523]), .out(
        \prgm_register/n1049 ) );
  nand2 \prgm_register/C4655  ( .a(\prgm_register/en_not ), .b(a[524]), .out(
        \prgm_register/n1050 ) );
  nand2 \prgm_register/C4656  ( .a(\prgm_register/n1049 ), .b(
        \prgm_register/n1050 ), .out(\prgm_register/or_signal [524]) );
  nand2 \prgm_register/C4657  ( .a(enable), .b(a[524]), .out(
        \prgm_register/n1051 ) );
  nand2 \prgm_register/C4658  ( .a(\prgm_register/en_not ), .b(a[525]), .out(
        \prgm_register/n1052 ) );
  nand2 \prgm_register/C4659  ( .a(\prgm_register/n1051 ), .b(
        \prgm_register/n1052 ), .out(\prgm_register/or_signal [525]) );
  nand2 \prgm_register/C4660  ( .a(enable), .b(a[525]), .out(
        \prgm_register/n1053 ) );
  nand2 \prgm_register/C4661  ( .a(\prgm_register/en_not ), .b(a[526]), .out(
        \prgm_register/n1054 ) );
  nand2 \prgm_register/C4662  ( .a(\prgm_register/n1053 ), .b(
        \prgm_register/n1054 ), .out(\prgm_register/or_signal [526]) );
  nand2 \prgm_register/C4663  ( .a(enable), .b(a[526]), .out(
        \prgm_register/n1055 ) );
  nand2 \prgm_register/C4664  ( .a(\prgm_register/en_not ), .b(a[527]), .out(
        \prgm_register/n1056 ) );
  nand2 \prgm_register/C4665  ( .a(\prgm_register/n1055 ), .b(
        \prgm_register/n1056 ), .out(\prgm_register/or_signal [527]) );
  nand2 \prgm_register/C4666  ( .a(enable), .b(a[527]), .out(
        \prgm_register/n1057 ) );
  nand2 \prgm_register/C4667  ( .a(\prgm_register/en_not ), .b(a[528]), .out(
        \prgm_register/n1058 ) );
  nand2 \prgm_register/C4668  ( .a(\prgm_register/n1057 ), .b(
        \prgm_register/n1058 ), .out(\prgm_register/or_signal [528]) );
  nand2 \prgm_register/C4669  ( .a(enable), .b(a[528]), .out(
        \prgm_register/n1059 ) );
  nand2 \prgm_register/C4670  ( .a(\prgm_register/en_not ), .b(a[529]), .out(
        \prgm_register/n1060 ) );
  nand2 \prgm_register/C4671  ( .a(\prgm_register/n1059 ), .b(
        \prgm_register/n1060 ), .out(\prgm_register/or_signal [529]) );
  nand2 \prgm_register/C4672  ( .a(enable), .b(a[529]), .out(
        \prgm_register/n1061 ) );
  nand2 \prgm_register/C4673  ( .a(\prgm_register/en_not ), .b(a[530]), .out(
        \prgm_register/n1062 ) );
  nand2 \prgm_register/C4674  ( .a(\prgm_register/n1061 ), .b(
        \prgm_register/n1062 ), .out(\prgm_register/or_signal [530]) );
  nand2 \prgm_register/C4675  ( .a(enable), .b(a[530]), .out(
        \prgm_register/n1063 ) );
  nand2 \prgm_register/C4676  ( .a(\prgm_register/en_not ), .b(a[531]), .out(
        \prgm_register/n1064 ) );
  nand2 \prgm_register/C4677  ( .a(\prgm_register/n1063 ), .b(
        \prgm_register/n1064 ), .out(\prgm_register/or_signal [531]) );
  nand2 \prgm_register/C4678  ( .a(enable), .b(a[531]), .out(
        \prgm_register/n1065 ) );
  nand2 \prgm_register/C4679  ( .a(\prgm_register/en_not ), .b(a[532]), .out(
        \prgm_register/n1066 ) );
  nand2 \prgm_register/C4680  ( .a(\prgm_register/n1065 ), .b(
        \prgm_register/n1066 ), .out(\prgm_register/or_signal [532]) );
  nand2 \prgm_register/C4681  ( .a(enable), .b(a[532]), .out(
        \prgm_register/n1067 ) );
  nand2 \prgm_register/C4682  ( .a(\prgm_register/en_not ), .b(a[533]), .out(
        \prgm_register/n1068 ) );
  nand2 \prgm_register/C4683  ( .a(\prgm_register/n1067 ), .b(
        \prgm_register/n1068 ), .out(\prgm_register/or_signal [533]) );
  nand2 \prgm_register/C4684  ( .a(enable), .b(a[533]), .out(
        \prgm_register/n1069 ) );
  nand2 \prgm_register/C4685  ( .a(\prgm_register/en_not ), .b(a[534]), .out(
        \prgm_register/n1070 ) );
  nand2 \prgm_register/C4686  ( .a(\prgm_register/n1069 ), .b(
        \prgm_register/n1070 ), .out(\prgm_register/or_signal [534]) );
  nand2 \prgm_register/C4687  ( .a(enable), .b(a[534]), .out(
        \prgm_register/n1071 ) );
  nand2 \prgm_register/C4688  ( .a(\prgm_register/en_not ), .b(a[535]), .out(
        \prgm_register/n1072 ) );
  nand2 \prgm_register/C4689  ( .a(\prgm_register/n1071 ), .b(
        \prgm_register/n1072 ), .out(\prgm_register/or_signal [535]) );
  nand2 \prgm_register/C4690  ( .a(enable), .b(a[535]), .out(
        \prgm_register/n1073 ) );
  nand2 \prgm_register/C4691  ( .a(\prgm_register/en_not ), .b(a[536]), .out(
        \prgm_register/n1074 ) );
  nand2 \prgm_register/C4692  ( .a(\prgm_register/n1073 ), .b(
        \prgm_register/n1074 ), .out(\prgm_register/or_signal [536]) );
  nand2 \prgm_register/C4693  ( .a(enable), .b(a[536]), .out(
        \prgm_register/n1075 ) );
  nand2 \prgm_register/C4694  ( .a(\prgm_register/en_not ), .b(a[537]), .out(
        \prgm_register/n1076 ) );
  nand2 \prgm_register/C4695  ( .a(\prgm_register/n1075 ), .b(
        \prgm_register/n1076 ), .out(\prgm_register/or_signal [537]) );
  nand2 \prgm_register/C4696  ( .a(enable), .b(a[537]), .out(
        \prgm_register/n1077 ) );
  nand2 \prgm_register/C4697  ( .a(\prgm_register/en_not ), .b(a[538]), .out(
        \prgm_register/n1078 ) );
  nand2 \prgm_register/C4698  ( .a(\prgm_register/n1077 ), .b(
        \prgm_register/n1078 ), .out(\prgm_register/or_signal [538]) );
  nand2 \prgm_register/C4699  ( .a(enable), .b(a[538]), .out(
        \prgm_register/n1079 ) );
  nand2 \prgm_register/C4700  ( .a(\prgm_register/en_not ), .b(a[539]), .out(
        \prgm_register/n1080 ) );
  nand2 \prgm_register/C4701  ( .a(\prgm_register/n1079 ), .b(
        \prgm_register/n1080 ), .out(\prgm_register/or_signal [539]) );
  nand2 \prgm_register/C4702  ( .a(enable), .b(a[539]), .out(
        \prgm_register/n1081 ) );
  nand2 \prgm_register/C4703  ( .a(\prgm_register/en_not ), .b(a[540]), .out(
        \prgm_register/n1082 ) );
  nand2 \prgm_register/C4704  ( .a(\prgm_register/n1081 ), .b(
        \prgm_register/n1082 ), .out(\prgm_register/or_signal [540]) );
  nand2 \prgm_register/C4705  ( .a(enable), .b(a[540]), .out(
        \prgm_register/n1083 ) );
  nand2 \prgm_register/C4706  ( .a(\prgm_register/en_not ), .b(a[541]), .out(
        \prgm_register/n1084 ) );
  nand2 \prgm_register/C4707  ( .a(\prgm_register/n1083 ), .b(
        \prgm_register/n1084 ), .out(\prgm_register/or_signal [541]) );
  nand2 \prgm_register/C4708  ( .a(enable), .b(a[541]), .out(
        \prgm_register/n1085 ) );
  nand2 \prgm_register/C4709  ( .a(\prgm_register/en_not ), .b(a[542]), .out(
        \prgm_register/n1086 ) );
  nand2 \prgm_register/C4710  ( .a(\prgm_register/n1085 ), .b(
        \prgm_register/n1086 ), .out(\prgm_register/or_signal [542]) );
  nand2 \prgm_register/C4711  ( .a(enable), .b(a[542]), .out(
        \prgm_register/n1087 ) );
  nand2 \prgm_register/C4712  ( .a(\prgm_register/en_not ), .b(a[543]), .out(
        \prgm_register/n1088 ) );
  nand2 \prgm_register/C4713  ( .a(\prgm_register/n1087 ), .b(
        \prgm_register/n1088 ), .out(\prgm_register/or_signal [543]) );
  nand2 \prgm_register/C4714  ( .a(enable), .b(a[543]), .out(
        \prgm_register/n1089 ) );
  nand2 \prgm_register/C4715  ( .a(\prgm_register/en_not ), .b(a[544]), .out(
        \prgm_register/n1090 ) );
  nand2 \prgm_register/C4716  ( .a(\prgm_register/n1089 ), .b(
        \prgm_register/n1090 ), .out(\prgm_register/or_signal [544]) );
  nand2 \prgm_register/C4717  ( .a(enable), .b(a[544]), .out(
        \prgm_register/n1091 ) );
  nand2 \prgm_register/C4718  ( .a(\prgm_register/en_not ), .b(a[545]), .out(
        \prgm_register/n1092 ) );
  nand2 \prgm_register/C4719  ( .a(\prgm_register/n1091 ), .b(
        \prgm_register/n1092 ), .out(\prgm_register/or_signal [545]) );
  nand2 \prgm_register/C4720  ( .a(enable), .b(a[545]), .out(
        \prgm_register/n1093 ) );
  nand2 \prgm_register/C4721  ( .a(\prgm_register/en_not ), .b(a[546]), .out(
        \prgm_register/n1094 ) );
  nand2 \prgm_register/C4722  ( .a(\prgm_register/n1093 ), .b(
        \prgm_register/n1094 ), .out(\prgm_register/or_signal [546]) );
  nand2 \prgm_register/C4723  ( .a(enable), .b(a[546]), .out(
        \prgm_register/n1095 ) );
  nand2 \prgm_register/C4724  ( .a(\prgm_register/en_not ), .b(a[547]), .out(
        \prgm_register/n1096 ) );
  nand2 \prgm_register/C4725  ( .a(\prgm_register/n1095 ), .b(
        \prgm_register/n1096 ), .out(\prgm_register/or_signal [547]) );
  nand2 \prgm_register/C4726  ( .a(enable), .b(a[547]), .out(
        \prgm_register/n1097 ) );
  nand2 \prgm_register/C4727  ( .a(\prgm_register/en_not ), .b(a[548]), .out(
        \prgm_register/n1098 ) );
  nand2 \prgm_register/C4728  ( .a(\prgm_register/n1097 ), .b(
        \prgm_register/n1098 ), .out(\prgm_register/or_signal [548]) );
  nand2 \prgm_register/C4729  ( .a(enable), .b(a[548]), .out(
        \prgm_register/n1099 ) );
  nand2 \prgm_register/C4730  ( .a(\prgm_register/en_not ), .b(a[549]), .out(
        \prgm_register/n1100 ) );
  nand2 \prgm_register/C4731  ( .a(\prgm_register/n1099 ), .b(
        \prgm_register/n1100 ), .out(\prgm_register/or_signal [549]) );
  nand2 \prgm_register/C4732  ( .a(enable), .b(a[549]), .out(
        \prgm_register/n1101 ) );
  nand2 \prgm_register/C4733  ( .a(\prgm_register/en_not ), .b(a[550]), .out(
        \prgm_register/n1102 ) );
  nand2 \prgm_register/C4734  ( .a(\prgm_register/n1101 ), .b(
        \prgm_register/n1102 ), .out(\prgm_register/or_signal [550]) );
  nand2 \prgm_register/C4735  ( .a(enable), .b(a[550]), .out(
        \prgm_register/n1103 ) );
  nand2 \prgm_register/C4736  ( .a(\prgm_register/en_not ), .b(a[551]), .out(
        \prgm_register/n1104 ) );
  nand2 \prgm_register/C4737  ( .a(\prgm_register/n1103 ), .b(
        \prgm_register/n1104 ), .out(\prgm_register/or_signal [551]) );
  nand2 \prgm_register/C4738  ( .a(enable), .b(a[551]), .out(
        \prgm_register/n1105 ) );
  nand2 \prgm_register/C4739  ( .a(\prgm_register/en_not ), .b(a[552]), .out(
        \prgm_register/n1106 ) );
  nand2 \prgm_register/C4740  ( .a(\prgm_register/n1105 ), .b(
        \prgm_register/n1106 ), .out(\prgm_register/or_signal [552]) );
  nand2 \prgm_register/C4741  ( .a(enable), .b(a[552]), .out(
        \prgm_register/n1107 ) );
  nand2 \prgm_register/C4742  ( .a(\prgm_register/en_not ), .b(a[553]), .out(
        \prgm_register/n1108 ) );
  nand2 \prgm_register/C4743  ( .a(\prgm_register/n1107 ), .b(
        \prgm_register/n1108 ), .out(\prgm_register/or_signal [553]) );
  nand2 \prgm_register/C4744  ( .a(enable), .b(a[553]), .out(
        \prgm_register/n1109 ) );
  nand2 \prgm_register/C4745  ( .a(\prgm_register/en_not ), .b(a[554]), .out(
        \prgm_register/n1110 ) );
  nand2 \prgm_register/C4746  ( .a(\prgm_register/n1109 ), .b(
        \prgm_register/n1110 ), .out(\prgm_register/or_signal [554]) );
  nand2 \prgm_register/C4747  ( .a(enable), .b(a[554]), .out(
        \prgm_register/n1111 ) );
  nand2 \prgm_register/C4748  ( .a(\prgm_register/en_not ), .b(a[555]), .out(
        \prgm_register/n1112 ) );
  nand2 \prgm_register/C4749  ( .a(\prgm_register/n1111 ), .b(
        \prgm_register/n1112 ), .out(\prgm_register/or_signal [555]) );
  nand2 \prgm_register/C4750  ( .a(enable), .b(a[555]), .out(
        \prgm_register/n1113 ) );
  nand2 \prgm_register/C4751  ( .a(\prgm_register/en_not ), .b(a[556]), .out(
        \prgm_register/n1114 ) );
  nand2 \prgm_register/C4752  ( .a(\prgm_register/n1113 ), .b(
        \prgm_register/n1114 ), .out(\prgm_register/or_signal [556]) );
  nand2 \prgm_register/C4753  ( .a(enable), .b(a[556]), .out(
        \prgm_register/n1115 ) );
  nand2 \prgm_register/C4754  ( .a(\prgm_register/en_not ), .b(a[557]), .out(
        \prgm_register/n1116 ) );
  nand2 \prgm_register/C4755  ( .a(\prgm_register/n1115 ), .b(
        \prgm_register/n1116 ), .out(\prgm_register/or_signal [557]) );
  nand2 \prgm_register/C4756  ( .a(enable), .b(a[557]), .out(
        \prgm_register/n1117 ) );
  nand2 \prgm_register/C4757  ( .a(\prgm_register/en_not ), .b(a[558]), .out(
        \prgm_register/n1118 ) );
  nand2 \prgm_register/C4758  ( .a(\prgm_register/n1117 ), .b(
        \prgm_register/n1118 ), .out(\prgm_register/or_signal [558]) );
  nand2 \prgm_register/C4759  ( .a(enable), .b(a[558]), .out(
        \prgm_register/n1119 ) );
  nand2 \prgm_register/C4760  ( .a(\prgm_register/en_not ), .b(a[559]), .out(
        \prgm_register/n1120 ) );
  nand2 \prgm_register/C4761  ( .a(\prgm_register/n1119 ), .b(
        \prgm_register/n1120 ), .out(\prgm_register/or_signal [559]) );
  nand2 \prgm_register/C4762  ( .a(enable), .b(a[559]), .out(
        \prgm_register/n1121 ) );
  nand2 \prgm_register/C4763  ( .a(\prgm_register/en_not ), .b(a[560]), .out(
        \prgm_register/n1122 ) );
  nand2 \prgm_register/C4764  ( .a(\prgm_register/n1121 ), .b(
        \prgm_register/n1122 ), .out(\prgm_register/or_signal [560]) );
  nand2 \prgm_register/C4765  ( .a(enable), .b(a[560]), .out(
        \prgm_register/n1123 ) );
  nand2 \prgm_register/C4766  ( .a(\prgm_register/en_not ), .b(a[561]), .out(
        \prgm_register/n1124 ) );
  nand2 \prgm_register/C4767  ( .a(\prgm_register/n1123 ), .b(
        \prgm_register/n1124 ), .out(\prgm_register/or_signal [561]) );
  nand2 \prgm_register/C4768  ( .a(enable), .b(a[561]), .out(
        \prgm_register/n1125 ) );
  nand2 \prgm_register/C4769  ( .a(\prgm_register/en_not ), .b(a[562]), .out(
        \prgm_register/n1126 ) );
  nand2 \prgm_register/C4770  ( .a(\prgm_register/n1125 ), .b(
        \prgm_register/n1126 ), .out(\prgm_register/or_signal [562]) );
  nand2 \prgm_register/C4771  ( .a(enable), .b(a[562]), .out(
        \prgm_register/n1127 ) );
  nand2 \prgm_register/C4772  ( .a(\prgm_register/en_not ), .b(a[563]), .out(
        \prgm_register/n1128 ) );
  nand2 \prgm_register/C4773  ( .a(\prgm_register/n1127 ), .b(
        \prgm_register/n1128 ), .out(\prgm_register/or_signal [563]) );
  nand2 \prgm_register/C4774  ( .a(enable), .b(a[563]), .out(
        \prgm_register/n1129 ) );
  nand2 \prgm_register/C4775  ( .a(\prgm_register/en_not ), .b(a[564]), .out(
        \prgm_register/n1130 ) );
  nand2 \prgm_register/C4776  ( .a(\prgm_register/n1129 ), .b(
        \prgm_register/n1130 ), .out(\prgm_register/or_signal [564]) );
  nand2 \prgm_register/C4777  ( .a(enable), .b(a[564]), .out(
        \prgm_register/n1131 ) );
  nand2 \prgm_register/C4778  ( .a(\prgm_register/en_not ), .b(a[565]), .out(
        \prgm_register/n1132 ) );
  nand2 \prgm_register/C4779  ( .a(\prgm_register/n1131 ), .b(
        \prgm_register/n1132 ), .out(\prgm_register/or_signal [565]) );
  nand2 \prgm_register/C4780  ( .a(enable), .b(a[565]), .out(
        \prgm_register/n1133 ) );
  nand2 \prgm_register/C4781  ( .a(\prgm_register/en_not ), .b(a[566]), .out(
        \prgm_register/n1134 ) );
  nand2 \prgm_register/C4782  ( .a(\prgm_register/n1133 ), .b(
        \prgm_register/n1134 ), .out(\prgm_register/or_signal [566]) );
  nand2 \prgm_register/C4783  ( .a(enable), .b(a[566]), .out(
        \prgm_register/n1135 ) );
  nand2 \prgm_register/C4784  ( .a(\prgm_register/en_not ), .b(a[567]), .out(
        \prgm_register/n1136 ) );
  nand2 \prgm_register/C4785  ( .a(\prgm_register/n1135 ), .b(
        \prgm_register/n1136 ), .out(\prgm_register/or_signal [567]) );
  nand2 \prgm_register/C4786  ( .a(enable), .b(a[567]), .out(
        \prgm_register/n1137 ) );
  nand2 \prgm_register/C4787  ( .a(\prgm_register/en_not ), .b(a[568]), .out(
        \prgm_register/n1138 ) );
  nand2 \prgm_register/C4788  ( .a(\prgm_register/n1137 ), .b(
        \prgm_register/n1138 ), .out(\prgm_register/or_signal [568]) );
  nand2 \prgm_register/C4789  ( .a(enable), .b(a[568]), .out(
        \prgm_register/n1139 ) );
  nand2 \prgm_register/C4790  ( .a(\prgm_register/en_not ), .b(a[569]), .out(
        \prgm_register/n1140 ) );
  nand2 \prgm_register/C4791  ( .a(\prgm_register/n1139 ), .b(
        \prgm_register/n1140 ), .out(\prgm_register/or_signal [569]) );
  nand2 \prgm_register/C4792  ( .a(enable), .b(a[569]), .out(
        \prgm_register/n1141 ) );
  nand2 \prgm_register/C4793  ( .a(\prgm_register/en_not ), .b(a[570]), .out(
        \prgm_register/n1142 ) );
  nand2 \prgm_register/C4794  ( .a(\prgm_register/n1141 ), .b(
        \prgm_register/n1142 ), .out(\prgm_register/or_signal [570]) );
  nand2 \prgm_register/C4795  ( .a(enable), .b(a[570]), .out(
        \prgm_register/n1143 ) );
  nand2 \prgm_register/C4796  ( .a(\prgm_register/en_not ), .b(a[571]), .out(
        \prgm_register/n1144 ) );
  nand2 \prgm_register/C4797  ( .a(\prgm_register/n1143 ), .b(
        \prgm_register/n1144 ), .out(\prgm_register/or_signal [571]) );
  nand2 \prgm_register/C4798  ( .a(enable), .b(a[571]), .out(
        \prgm_register/n1145 ) );
  nand2 \prgm_register/C4799  ( .a(\prgm_register/en_not ), .b(a[572]), .out(
        \prgm_register/n1146 ) );
  nand2 \prgm_register/C4800  ( .a(\prgm_register/n1145 ), .b(
        \prgm_register/n1146 ), .out(\prgm_register/or_signal [572]) );
  nand2 \prgm_register/C4801  ( .a(enable), .b(a[572]), .out(
        \prgm_register/n1147 ) );
  nand2 \prgm_register/C4802  ( .a(\prgm_register/en_not ), .b(a[573]), .out(
        \prgm_register/n1148 ) );
  nand2 \prgm_register/C4803  ( .a(\prgm_register/n1147 ), .b(
        \prgm_register/n1148 ), .out(\prgm_register/or_signal [573]) );
  nand2 \prgm_register/C4804  ( .a(enable), .b(a[573]), .out(
        \prgm_register/n1149 ) );
  nand2 \prgm_register/C4805  ( .a(\prgm_register/en_not ), .b(a[574]), .out(
        \prgm_register/n1150 ) );
  nand2 \prgm_register/C4806  ( .a(\prgm_register/n1149 ), .b(
        \prgm_register/n1150 ), .out(\prgm_register/or_signal [574]) );
  nand2 \prgm_register/C4807  ( .a(enable), .b(a[574]), .out(
        \prgm_register/n1151 ) );
  nand2 \prgm_register/C4808  ( .a(\prgm_register/en_not ), .b(a[575]), .out(
        \prgm_register/n1152 ) );
  nand2 \prgm_register/C4809  ( .a(\prgm_register/n1151 ), .b(
        \prgm_register/n1152 ), .out(\prgm_register/or_signal [575]) );
  nand2 \prgm_register/C4810  ( .a(enable), .b(a[575]), .out(
        \prgm_register/n1153 ) );
  nand2 \prgm_register/C4811  ( .a(\prgm_register/en_not ), .b(a[576]), .out(
        \prgm_register/n1154 ) );
  nand2 \prgm_register/C4812  ( .a(\prgm_register/n1153 ), .b(
        \prgm_register/n1154 ), .out(\prgm_register/or_signal [576]) );
  nand2 \prgm_register/C4813  ( .a(enable), .b(a[576]), .out(
        \prgm_register/n1155 ) );
  nand2 \prgm_register/C4814  ( .a(\prgm_register/en_not ), .b(a[577]), .out(
        \prgm_register/n1156 ) );
  nand2 \prgm_register/C4815  ( .a(\prgm_register/n1155 ), .b(
        \prgm_register/n1156 ), .out(\prgm_register/or_signal [577]) );
  nand2 \prgm_register/C4816  ( .a(enable), .b(a[577]), .out(
        \prgm_register/n1157 ) );
  nand2 \prgm_register/C4817  ( .a(\prgm_register/en_not ), .b(a[578]), .out(
        \prgm_register/n1158 ) );
  nand2 \prgm_register/C4818  ( .a(\prgm_register/n1157 ), .b(
        \prgm_register/n1158 ), .out(\prgm_register/or_signal [578]) );
  nand2 \prgm_register/C4819  ( .a(enable), .b(a[578]), .out(
        \prgm_register/n1159 ) );
  nand2 \prgm_register/C4820  ( .a(\prgm_register/en_not ), .b(a[579]), .out(
        \prgm_register/n1160 ) );
  nand2 \prgm_register/C4821  ( .a(\prgm_register/n1159 ), .b(
        \prgm_register/n1160 ), .out(\prgm_register/or_signal [579]) );
  nand2 \prgm_register/C4822  ( .a(enable), .b(a[579]), .out(
        \prgm_register/n1161 ) );
  nand2 \prgm_register/C4823  ( .a(\prgm_register/en_not ), .b(a[580]), .out(
        \prgm_register/n1162 ) );
  nand2 \prgm_register/C4824  ( .a(\prgm_register/n1161 ), .b(
        \prgm_register/n1162 ), .out(\prgm_register/or_signal [580]) );
  nand2 \prgm_register/C4825  ( .a(enable), .b(a[580]), .out(
        \prgm_register/n1163 ) );
  nand2 \prgm_register/C4826  ( .a(\prgm_register/en_not ), .b(a[581]), .out(
        \prgm_register/n1164 ) );
  nand2 \prgm_register/C4827  ( .a(\prgm_register/n1163 ), .b(
        \prgm_register/n1164 ), .out(\prgm_register/or_signal [581]) );
  nand2 \prgm_register/C4828  ( .a(enable), .b(a[581]), .out(
        \prgm_register/n1165 ) );
  nand2 \prgm_register/C4829  ( .a(\prgm_register/en_not ), .b(a[582]), .out(
        \prgm_register/n1166 ) );
  nand2 \prgm_register/C4830  ( .a(\prgm_register/n1165 ), .b(
        \prgm_register/n1166 ), .out(\prgm_register/or_signal [582]) );
  nand2 \prgm_register/C4831  ( .a(enable), .b(a[582]), .out(
        \prgm_register/n1167 ) );
  nand2 \prgm_register/C4832  ( .a(\prgm_register/en_not ), .b(a[583]), .out(
        \prgm_register/n1168 ) );
  nand2 \prgm_register/C4833  ( .a(\prgm_register/n1167 ), .b(
        \prgm_register/n1168 ), .out(\prgm_register/or_signal [583]) );
  nand2 \prgm_register/C4834  ( .a(enable), .b(a[583]), .out(
        \prgm_register/n1169 ) );
  nand2 \prgm_register/C4835  ( .a(\prgm_register/en_not ), .b(a[584]), .out(
        \prgm_register/n1170 ) );
  nand2 \prgm_register/C4836  ( .a(\prgm_register/n1169 ), .b(
        \prgm_register/n1170 ), .out(\prgm_register/or_signal [584]) );
  nand2 \prgm_register/C4837  ( .a(enable), .b(a[584]), .out(
        \prgm_register/n1171 ) );
  nand2 \prgm_register/C4838  ( .a(\prgm_register/en_not ), .b(a[585]), .out(
        \prgm_register/n1172 ) );
  nand2 \prgm_register/C4839  ( .a(\prgm_register/n1171 ), .b(
        \prgm_register/n1172 ), .out(\prgm_register/or_signal [585]) );
  nand2 \prgm_register/C4840  ( .a(enable), .b(a[585]), .out(
        \prgm_register/n1173 ) );
  nand2 \prgm_register/C4841  ( .a(\prgm_register/en_not ), .b(a[586]), .out(
        \prgm_register/n1174 ) );
  nand2 \prgm_register/C4842  ( .a(\prgm_register/n1173 ), .b(
        \prgm_register/n1174 ), .out(\prgm_register/or_signal [586]) );
  nand2 \prgm_register/C4843  ( .a(enable), .b(a[586]), .out(
        \prgm_register/n1175 ) );
  nand2 \prgm_register/C4844  ( .a(\prgm_register/en_not ), .b(a[587]), .out(
        \prgm_register/n1176 ) );
  nand2 \prgm_register/C4845  ( .a(\prgm_register/n1175 ), .b(
        \prgm_register/n1176 ), .out(\prgm_register/or_signal [587]) );
  nand2 \prgm_register/C4846  ( .a(enable), .b(a[587]), .out(
        \prgm_register/n1177 ) );
  nand2 \prgm_register/C4847  ( .a(\prgm_register/en_not ), .b(a[588]), .out(
        \prgm_register/n1178 ) );
  nand2 \prgm_register/C4848  ( .a(\prgm_register/n1177 ), .b(
        \prgm_register/n1178 ), .out(\prgm_register/or_signal [588]) );
  nand2 \prgm_register/C4849  ( .a(enable), .b(a[588]), .out(
        \prgm_register/n1179 ) );
  nand2 \prgm_register/C4850  ( .a(\prgm_register/en_not ), .b(a[589]), .out(
        \prgm_register/n1180 ) );
  nand2 \prgm_register/C4851  ( .a(\prgm_register/n1179 ), .b(
        \prgm_register/n1180 ), .out(\prgm_register/or_signal [589]) );
  nand2 \prgm_register/C4852  ( .a(enable), .b(a[589]), .out(
        \prgm_register/n1181 ) );
  nand2 \prgm_register/C4853  ( .a(\prgm_register/en_not ), .b(a[590]), .out(
        \prgm_register/n1182 ) );
  nand2 \prgm_register/C4854  ( .a(\prgm_register/n1181 ), .b(
        \prgm_register/n1182 ), .out(\prgm_register/or_signal [590]) );
  nand2 \prgm_register/C4855  ( .a(enable), .b(a[590]), .out(
        \prgm_register/n1183 ) );
  nand2 \prgm_register/C4856  ( .a(\prgm_register/en_not ), .b(a[591]), .out(
        \prgm_register/n1184 ) );
  nand2 \prgm_register/C4857  ( .a(\prgm_register/n1183 ), .b(
        \prgm_register/n1184 ), .out(\prgm_register/or_signal [591]) );
  nand2 \prgm_register/C4858  ( .a(enable), .b(a[591]), .out(
        \prgm_register/n1185 ) );
  nand2 \prgm_register/C4859  ( .a(\prgm_register/en_not ), .b(a[592]), .out(
        \prgm_register/n1186 ) );
  nand2 \prgm_register/C4860  ( .a(\prgm_register/n1185 ), .b(
        \prgm_register/n1186 ), .out(\prgm_register/or_signal [592]) );
  nand2 \prgm_register/C4861  ( .a(enable), .b(a[592]), .out(
        \prgm_register/n1187 ) );
  nand2 \prgm_register/C4862  ( .a(\prgm_register/en_not ), .b(a[593]), .out(
        \prgm_register/n1188 ) );
  nand2 \prgm_register/C4863  ( .a(\prgm_register/n1187 ), .b(
        \prgm_register/n1188 ), .out(\prgm_register/or_signal [593]) );
  nand2 \prgm_register/C4864  ( .a(enable), .b(a[593]), .out(
        \prgm_register/n1189 ) );
  nand2 \prgm_register/C4865  ( .a(\prgm_register/en_not ), .b(a[594]), .out(
        \prgm_register/n1190 ) );
  nand2 \prgm_register/C4866  ( .a(\prgm_register/n1189 ), .b(
        \prgm_register/n1190 ), .out(\prgm_register/or_signal [594]) );
  nand2 \prgm_register/C4867  ( .a(enable), .b(a[594]), .out(
        \prgm_register/n1191 ) );
  nand2 \prgm_register/C4868  ( .a(\prgm_register/en_not ), .b(a[595]), .out(
        \prgm_register/n1192 ) );
  nand2 \prgm_register/C4869  ( .a(\prgm_register/n1191 ), .b(
        \prgm_register/n1192 ), .out(\prgm_register/or_signal [595]) );
  nand2 \prgm_register/C4870  ( .a(enable), .b(a[595]), .out(
        \prgm_register/n1193 ) );
  nand2 \prgm_register/C4871  ( .a(\prgm_register/en_not ), .b(a[596]), .out(
        \prgm_register/n1194 ) );
  nand2 \prgm_register/C4872  ( .a(\prgm_register/n1193 ), .b(
        \prgm_register/n1194 ), .out(\prgm_register/or_signal [596]) );
  nand2 \prgm_register/C4873  ( .a(enable), .b(a[596]), .out(
        \prgm_register/n1195 ) );
  nand2 \prgm_register/C4874  ( .a(\prgm_register/en_not ), .b(a[597]), .out(
        \prgm_register/n1196 ) );
  nand2 \prgm_register/C4875  ( .a(\prgm_register/n1195 ), .b(
        \prgm_register/n1196 ), .out(\prgm_register/or_signal [597]) );
  nand2 \prgm_register/C4876  ( .a(enable), .b(a[597]), .out(
        \prgm_register/n1197 ) );
  nand2 \prgm_register/C4877  ( .a(\prgm_register/en_not ), .b(a[598]), .out(
        \prgm_register/n1198 ) );
  nand2 \prgm_register/C4878  ( .a(\prgm_register/n1197 ), .b(
        \prgm_register/n1198 ), .out(\prgm_register/or_signal [598]) );
  nand2 \prgm_register/C4879  ( .a(enable), .b(a[598]), .out(
        \prgm_register/n1199 ) );
  nand2 \prgm_register/C4880  ( .a(\prgm_register/en_not ), .b(a[599]), .out(
        \prgm_register/n1200 ) );
  nand2 \prgm_register/C4881  ( .a(\prgm_register/n1199 ), .b(
        \prgm_register/n1200 ), .out(\prgm_register/or_signal [599]) );
  nand2 \prgm_register/C4882  ( .a(enable), .b(a[599]), .out(
        \prgm_register/n1201 ) );
  nand2 \prgm_register/C4883  ( .a(\prgm_register/en_not ), .b(a[600]), .out(
        \prgm_register/n1202 ) );
  nand2 \prgm_register/C4884  ( .a(\prgm_register/n1201 ), .b(
        \prgm_register/n1202 ), .out(\prgm_register/or_signal [600]) );
  nand2 \prgm_register/C4885  ( .a(enable), .b(a[600]), .out(
        \prgm_register/n1203 ) );
  nand2 \prgm_register/C4886  ( .a(\prgm_register/en_not ), .b(a[601]), .out(
        \prgm_register/n1204 ) );
  nand2 \prgm_register/C4887  ( .a(\prgm_register/n1203 ), .b(
        \prgm_register/n1204 ), .out(\prgm_register/or_signal [601]) );
  nand2 \prgm_register/C4888  ( .a(enable), .b(a[601]), .out(
        \prgm_register/n1205 ) );
  nand2 \prgm_register/C4889  ( .a(\prgm_register/en_not ), .b(a[602]), .out(
        \prgm_register/n1206 ) );
  nand2 \prgm_register/C4890  ( .a(\prgm_register/n1205 ), .b(
        \prgm_register/n1206 ), .out(\prgm_register/or_signal [602]) );
  nand2 \prgm_register/C4891  ( .a(enable), .b(a[602]), .out(
        \prgm_register/n1207 ) );
  nand2 \prgm_register/C4892  ( .a(\prgm_register/en_not ), .b(a[603]), .out(
        \prgm_register/n1208 ) );
  nand2 \prgm_register/C4893  ( .a(\prgm_register/n1207 ), .b(
        \prgm_register/n1208 ), .out(\prgm_register/or_signal [603]) );
  nand2 \prgm_register/C4894  ( .a(enable), .b(a[603]), .out(
        \prgm_register/n1209 ) );
  nand2 \prgm_register/C4895  ( .a(\prgm_register/en_not ), .b(a[604]), .out(
        \prgm_register/n1210 ) );
  nand2 \prgm_register/C4896  ( .a(\prgm_register/n1209 ), .b(
        \prgm_register/n1210 ), .out(\prgm_register/or_signal [604]) );
  nand2 \prgm_register/C4897  ( .a(enable), .b(a[604]), .out(
        \prgm_register/n1211 ) );
  nand2 \prgm_register/C4898  ( .a(\prgm_register/en_not ), .b(a[605]), .out(
        \prgm_register/n1212 ) );
  nand2 \prgm_register/C4899  ( .a(\prgm_register/n1211 ), .b(
        \prgm_register/n1212 ), .out(\prgm_register/or_signal [605]) );
  nand2 \prgm_register/C4900  ( .a(enable), .b(a[605]), .out(
        \prgm_register/n1213 ) );
  nand2 \prgm_register/C4901  ( .a(\prgm_register/en_not ), .b(a[606]), .out(
        \prgm_register/n1214 ) );
  nand2 \prgm_register/C4902  ( .a(\prgm_register/n1213 ), .b(
        \prgm_register/n1214 ), .out(\prgm_register/or_signal [606]) );
  nand2 \prgm_register/C4903  ( .a(enable), .b(a[606]), .out(
        \prgm_register/n1215 ) );
  nand2 \prgm_register/C4904  ( .a(\prgm_register/en_not ), .b(a[607]), .out(
        \prgm_register/n1216 ) );
  nand2 \prgm_register/C4905  ( .a(\prgm_register/n1215 ), .b(
        \prgm_register/n1216 ), .out(\prgm_register/or_signal [607]) );
  nand2 \prgm_register/C4906  ( .a(enable), .b(a[607]), .out(
        \prgm_register/n1217 ) );
  nand2 \prgm_register/C4907  ( .a(\prgm_register/en_not ), .b(a[608]), .out(
        \prgm_register/n1218 ) );
  nand2 \prgm_register/C4908  ( .a(\prgm_register/n1217 ), .b(
        \prgm_register/n1218 ), .out(\prgm_register/or_signal [608]) );
  nand2 \prgm_register/C4909  ( .a(enable), .b(a[608]), .out(
        \prgm_register/n1219 ) );
  nand2 \prgm_register/C4910  ( .a(\prgm_register/en_not ), .b(a[609]), .out(
        \prgm_register/n1220 ) );
  nand2 \prgm_register/C4911  ( .a(\prgm_register/n1219 ), .b(
        \prgm_register/n1220 ), .out(\prgm_register/or_signal [609]) );
  nand2 \prgm_register/C4912  ( .a(enable), .b(a[609]), .out(
        \prgm_register/n1221 ) );
  nand2 \prgm_register/C4913  ( .a(\prgm_register/en_not ), .b(a[610]), .out(
        \prgm_register/n1222 ) );
  nand2 \prgm_register/C4914  ( .a(\prgm_register/n1221 ), .b(
        \prgm_register/n1222 ), .out(\prgm_register/or_signal [610]) );
  nand2 \prgm_register/C4915  ( .a(enable), .b(a[610]), .out(
        \prgm_register/n1223 ) );
  nand2 \prgm_register/C4916  ( .a(\prgm_register/en_not ), .b(a[611]), .out(
        \prgm_register/n1224 ) );
  nand2 \prgm_register/C4917  ( .a(\prgm_register/n1223 ), .b(
        \prgm_register/n1224 ), .out(\prgm_register/or_signal [611]) );
  nand2 \prgm_register/C4918  ( .a(enable), .b(a[611]), .out(
        \prgm_register/n1225 ) );
  nand2 \prgm_register/C4919  ( .a(\prgm_register/en_not ), .b(a[612]), .out(
        \prgm_register/n1226 ) );
  nand2 \prgm_register/C4920  ( .a(\prgm_register/n1225 ), .b(
        \prgm_register/n1226 ), .out(\prgm_register/or_signal [612]) );
  nand2 \prgm_register/C4921  ( .a(enable), .b(a[612]), .out(
        \prgm_register/n1227 ) );
  nand2 \prgm_register/C4922  ( .a(\prgm_register/en_not ), .b(a[613]), .out(
        \prgm_register/n1228 ) );
  nand2 \prgm_register/C4923  ( .a(\prgm_register/n1227 ), .b(
        \prgm_register/n1228 ), .out(\prgm_register/or_signal [613]) );
  nand2 \prgm_register/C4924  ( .a(enable), .b(a[613]), .out(
        \prgm_register/n1229 ) );
  nand2 \prgm_register/C4925  ( .a(\prgm_register/en_not ), .b(a[614]), .out(
        \prgm_register/n1230 ) );
  nand2 \prgm_register/C4926  ( .a(\prgm_register/n1229 ), .b(
        \prgm_register/n1230 ), .out(\prgm_register/or_signal [614]) );
  nand2 \prgm_register/C4927  ( .a(enable), .b(a[614]), .out(
        \prgm_register/n1231 ) );
  nand2 \prgm_register/C4928  ( .a(\prgm_register/en_not ), .b(a[615]), .out(
        \prgm_register/n1232 ) );
  nand2 \prgm_register/C4929  ( .a(\prgm_register/n1231 ), .b(
        \prgm_register/n1232 ), .out(\prgm_register/or_signal [615]) );
  nand2 \prgm_register/C4930  ( .a(enable), .b(a[615]), .out(
        \prgm_register/n1233 ) );
  nand2 \prgm_register/C4931  ( .a(\prgm_register/en_not ), .b(a[616]), .out(
        \prgm_register/n1234 ) );
  nand2 \prgm_register/C4932  ( .a(\prgm_register/n1233 ), .b(
        \prgm_register/n1234 ), .out(\prgm_register/or_signal [616]) );
  nand2 \prgm_register/C4933  ( .a(enable), .b(a[616]), .out(
        \prgm_register/n1235 ) );
  nand2 \prgm_register/C4934  ( .a(\prgm_register/en_not ), .b(a[617]), .out(
        \prgm_register/n1236 ) );
  nand2 \prgm_register/C4935  ( .a(\prgm_register/n1235 ), .b(
        \prgm_register/n1236 ), .out(\prgm_register/or_signal [617]) );
  nand2 \prgm_register/C4936  ( .a(enable), .b(a[617]), .out(
        \prgm_register/n1237 ) );
  nand2 \prgm_register/C4937  ( .a(\prgm_register/en_not ), .b(a[618]), .out(
        \prgm_register/n1238 ) );
  nand2 \prgm_register/C4938  ( .a(\prgm_register/n1237 ), .b(
        \prgm_register/n1238 ), .out(\prgm_register/or_signal [618]) );
  nand2 \prgm_register/C4939  ( .a(enable), .b(a[618]), .out(
        \prgm_register/n1239 ) );
  nand2 \prgm_register/C4940  ( .a(\prgm_register/en_not ), .b(a[619]), .out(
        \prgm_register/n1240 ) );
  nand2 \prgm_register/C4941  ( .a(\prgm_register/n1239 ), .b(
        \prgm_register/n1240 ), .out(\prgm_register/or_signal [619]) );
  nand2 \prgm_register/C4942  ( .a(enable), .b(a[619]), .out(
        \prgm_register/n1241 ) );
  nand2 \prgm_register/C4943  ( .a(\prgm_register/en_not ), .b(a[620]), .out(
        \prgm_register/n1242 ) );
  nand2 \prgm_register/C4944  ( .a(\prgm_register/n1241 ), .b(
        \prgm_register/n1242 ), .out(\prgm_register/or_signal [620]) );
  nand2 \prgm_register/C4945  ( .a(enable), .b(a[620]), .out(
        \prgm_register/n1243 ) );
  nand2 \prgm_register/C4946  ( .a(\prgm_register/en_not ), .b(a[621]), .out(
        \prgm_register/n1244 ) );
  nand2 \prgm_register/C4947  ( .a(\prgm_register/n1243 ), .b(
        \prgm_register/n1244 ), .out(\prgm_register/or_signal [621]) );
  nand2 \prgm_register/C4948  ( .a(enable), .b(a[621]), .out(
        \prgm_register/n1245 ) );
  nand2 \prgm_register/C4949  ( .a(\prgm_register/en_not ), .b(a[622]), .out(
        \prgm_register/n1246 ) );
  nand2 \prgm_register/C4950  ( .a(\prgm_register/n1245 ), .b(
        \prgm_register/n1246 ), .out(\prgm_register/or_signal [622]) );
  nand2 \prgm_register/C4951  ( .a(enable), .b(a[622]), .out(
        \prgm_register/n1247 ) );
  nand2 \prgm_register/C4952  ( .a(\prgm_register/en_not ), .b(a[623]), .out(
        \prgm_register/n1248 ) );
  nand2 \prgm_register/C4953  ( .a(\prgm_register/n1247 ), .b(
        \prgm_register/n1248 ), .out(\prgm_register/or_signal [623]) );
  nand2 \prgm_register/C4954  ( .a(enable), .b(a[623]), .out(
        \prgm_register/n1249 ) );
  nand2 \prgm_register/C4955  ( .a(\prgm_register/en_not ), .b(a[624]), .out(
        \prgm_register/n1250 ) );
  nand2 \prgm_register/C4956  ( .a(\prgm_register/n1249 ), .b(
        \prgm_register/n1250 ), .out(\prgm_register/or_signal [624]) );
  nand2 \prgm_register/C4957  ( .a(enable), .b(a[624]), .out(
        \prgm_register/n1251 ) );
  nand2 \prgm_register/C4958  ( .a(\prgm_register/en_not ), .b(a[625]), .out(
        \prgm_register/n1252 ) );
  nand2 \prgm_register/C4959  ( .a(\prgm_register/n1251 ), .b(
        \prgm_register/n1252 ), .out(\prgm_register/or_signal [625]) );
  nand2 \prgm_register/C4960  ( .a(enable), .b(a[625]), .out(
        \prgm_register/n1253 ) );
  nand2 \prgm_register/C4961  ( .a(\prgm_register/en_not ), .b(a[626]), .out(
        \prgm_register/n1254 ) );
  nand2 \prgm_register/C4962  ( .a(\prgm_register/n1253 ), .b(
        \prgm_register/n1254 ), .out(\prgm_register/or_signal [626]) );
  nand2 \prgm_register/C4963  ( .a(enable), .b(a[626]), .out(
        \prgm_register/n1255 ) );
  nand2 \prgm_register/C4964  ( .a(\prgm_register/en_not ), .b(a[627]), .out(
        \prgm_register/n1256 ) );
  nand2 \prgm_register/C4965  ( .a(\prgm_register/n1255 ), .b(
        \prgm_register/n1256 ), .out(\prgm_register/or_signal [627]) );
  nand2 \prgm_register/C4966  ( .a(enable), .b(a[627]), .out(
        \prgm_register/n1257 ) );
  nand2 \prgm_register/C4967  ( .a(\prgm_register/en_not ), .b(a[628]), .out(
        \prgm_register/n1258 ) );
  nand2 \prgm_register/C4968  ( .a(\prgm_register/n1257 ), .b(
        \prgm_register/n1258 ), .out(\prgm_register/or_signal [628]) );
  nand2 \prgm_register/C4969  ( .a(enable), .b(a[628]), .out(
        \prgm_register/n1259 ) );
  nand2 \prgm_register/C4970  ( .a(\prgm_register/en_not ), .b(a[629]), .out(
        \prgm_register/n1260 ) );
  nand2 \prgm_register/C4971  ( .a(\prgm_register/n1259 ), .b(
        \prgm_register/n1260 ), .out(\prgm_register/or_signal [629]) );
  nand2 \prgm_register/C4972  ( .a(enable), .b(a[629]), .out(
        \prgm_register/n1261 ) );
  nand2 \prgm_register/C4973  ( .a(\prgm_register/en_not ), .b(a[630]), .out(
        \prgm_register/n1262 ) );
  nand2 \prgm_register/C4974  ( .a(\prgm_register/n1261 ), .b(
        \prgm_register/n1262 ), .out(\prgm_register/or_signal [630]) );
  nand2 \prgm_register/C4975  ( .a(enable), .b(a[630]), .out(
        \prgm_register/n1263 ) );
  nand2 \prgm_register/C4976  ( .a(\prgm_register/en_not ), .b(a[631]), .out(
        \prgm_register/n1264 ) );
  nand2 \prgm_register/C4977  ( .a(\prgm_register/n1263 ), .b(
        \prgm_register/n1264 ), .out(\prgm_register/or_signal [631]) );
  nand2 \prgm_register/C4978  ( .a(enable), .b(a[631]), .out(
        \prgm_register/n1265 ) );
  nand2 \prgm_register/C4979  ( .a(\prgm_register/en_not ), .b(a[632]), .out(
        \prgm_register/n1266 ) );
  nand2 \prgm_register/C4980  ( .a(\prgm_register/n1265 ), .b(
        \prgm_register/n1266 ), .out(\prgm_register/or_signal [632]) );
  nand2 \prgm_register/C4981  ( .a(enable), .b(a[632]), .out(
        \prgm_register/n1267 ) );
  nand2 \prgm_register/C4982  ( .a(\prgm_register/en_not ), .b(a[633]), .out(
        \prgm_register/n1268 ) );
  nand2 \prgm_register/C4983  ( .a(\prgm_register/n1267 ), .b(
        \prgm_register/n1268 ), .out(\prgm_register/or_signal [633]) );
  nand2 \prgm_register/C4984  ( .a(enable), .b(a[633]), .out(
        \prgm_register/n1269 ) );
  nand2 \prgm_register/C4985  ( .a(\prgm_register/en_not ), .b(a[634]), .out(
        \prgm_register/n1270 ) );
  nand2 \prgm_register/C4986  ( .a(\prgm_register/n1269 ), .b(
        \prgm_register/n1270 ), .out(\prgm_register/or_signal [634]) );
  nand2 \prgm_register/C4987  ( .a(enable), .b(a[634]), .out(
        \prgm_register/n1271 ) );
  nand2 \prgm_register/C4988  ( .a(\prgm_register/en_not ), .b(a[635]), .out(
        \prgm_register/n1272 ) );
  nand2 \prgm_register/C4989  ( .a(\prgm_register/n1271 ), .b(
        \prgm_register/n1272 ), .out(\prgm_register/or_signal [635]) );
  nand2 \prgm_register/C4990  ( .a(enable), .b(a[635]), .out(
        \prgm_register/n1273 ) );
  nand2 \prgm_register/C4991  ( .a(\prgm_register/en_not ), .b(a[636]), .out(
        \prgm_register/n1274 ) );
  nand2 \prgm_register/C4992  ( .a(\prgm_register/n1273 ), .b(
        \prgm_register/n1274 ), .out(\prgm_register/or_signal [636]) );
  nand2 \prgm_register/C4993  ( .a(enable), .b(a[636]), .out(
        \prgm_register/n1275 ) );
  nand2 \prgm_register/C4994  ( .a(\prgm_register/en_not ), .b(a[637]), .out(
        \prgm_register/n1276 ) );
  nand2 \prgm_register/C4995  ( .a(\prgm_register/n1275 ), .b(
        \prgm_register/n1276 ), .out(\prgm_register/or_signal [637]) );
  nand2 \prgm_register/C4996  ( .a(enable), .b(a[637]), .out(
        \prgm_register/n1277 ) );
  nand2 \prgm_register/C4997  ( .a(\prgm_register/en_not ), .b(a[638]), .out(
        \prgm_register/n1278 ) );
  nand2 \prgm_register/C4998  ( .a(\prgm_register/n1277 ), .b(
        \prgm_register/n1278 ), .out(\prgm_register/or_signal [638]) );
  nand2 \prgm_register/C4999  ( .a(enable), .b(a[638]), .out(
        \prgm_register/n1279 ) );
  nand2 \prgm_register/C5000  ( .a(\prgm_register/en_not ), .b(a[639]), .out(
        \prgm_register/n1280 ) );
  nand2 \prgm_register/C5001  ( .a(\prgm_register/n1279 ), .b(
        \prgm_register/n1280 ), .out(\prgm_register/or_signal [639]) );
  nand2 \prgm_register/C5002  ( .a(enable), .b(a[639]), .out(
        \prgm_register/n1281 ) );
  nand2 \prgm_register/C5003  ( .a(\prgm_register/en_not ), .b(a[640]), .out(
        \prgm_register/n1282 ) );
  nand2 \prgm_register/C5004  ( .a(\prgm_register/n1281 ), .b(
        \prgm_register/n1282 ), .out(\prgm_register/or_signal [640]) );
  nand2 \prgm_register/C5005  ( .a(enable), .b(a[640]), .out(
        \prgm_register/n1283 ) );
  nand2 \prgm_register/C5006  ( .a(\prgm_register/en_not ), .b(a[641]), .out(
        \prgm_register/n1284 ) );
  nand2 \prgm_register/C5007  ( .a(\prgm_register/n1283 ), .b(
        \prgm_register/n1284 ), .out(\prgm_register/or_signal [641]) );
  nand2 \prgm_register/C5008  ( .a(enable), .b(a[641]), .out(
        \prgm_register/n1285 ) );
  nand2 \prgm_register/C5009  ( .a(\prgm_register/en_not ), .b(a[642]), .out(
        \prgm_register/n1286 ) );
  nand2 \prgm_register/C5010  ( .a(\prgm_register/n1285 ), .b(
        \prgm_register/n1286 ), .out(\prgm_register/or_signal [642]) );
  nand2 \prgm_register/C5011  ( .a(enable), .b(a[642]), .out(
        \prgm_register/n1287 ) );
  nand2 \prgm_register/C5012  ( .a(\prgm_register/en_not ), .b(a[643]), .out(
        \prgm_register/n1288 ) );
  nand2 \prgm_register/C5013  ( .a(\prgm_register/n1287 ), .b(
        \prgm_register/n1288 ), .out(\prgm_register/or_signal [643]) );
  nand2 \prgm_register/C5014  ( .a(enable), .b(a[643]), .out(
        \prgm_register/n1289 ) );
  nand2 \prgm_register/C5015  ( .a(\prgm_register/en_not ), .b(a[644]), .out(
        \prgm_register/n1290 ) );
  nand2 \prgm_register/C5016  ( .a(\prgm_register/n1289 ), .b(
        \prgm_register/n1290 ), .out(\prgm_register/or_signal [644]) );
  nand2 \prgm_register/C5017  ( .a(enable), .b(a[644]), .out(
        \prgm_register/n1291 ) );
  nand2 \prgm_register/C5018  ( .a(\prgm_register/en_not ), .b(a[645]), .out(
        \prgm_register/n1292 ) );
  nand2 \prgm_register/C5019  ( .a(\prgm_register/n1291 ), .b(
        \prgm_register/n1292 ), .out(\prgm_register/or_signal [645]) );
  nand2 \prgm_register/C5020  ( .a(enable), .b(a[645]), .out(
        \prgm_register/n1293 ) );
  nand2 \prgm_register/C5021  ( .a(\prgm_register/en_not ), .b(a[646]), .out(
        \prgm_register/n1294 ) );
  nand2 \prgm_register/C5022  ( .a(\prgm_register/n1293 ), .b(
        \prgm_register/n1294 ), .out(\prgm_register/or_signal [646]) );
  nand2 \prgm_register/C5023  ( .a(enable), .b(a[646]), .out(
        \prgm_register/n1295 ) );
  nand2 \prgm_register/C5024  ( .a(\prgm_register/en_not ), .b(a[647]), .out(
        \prgm_register/n1296 ) );
  nand2 \prgm_register/C5025  ( .a(\prgm_register/n1295 ), .b(
        \prgm_register/n1296 ), .out(\prgm_register/or_signal [647]) );
  nand2 \prgm_register/C5026  ( .a(enable), .b(a[647]), .out(
        \prgm_register/n1297 ) );
  nand2 \prgm_register/C5027  ( .a(\prgm_register/en_not ), .b(a[648]), .out(
        \prgm_register/n1298 ) );
  nand2 \prgm_register/C5028  ( .a(\prgm_register/n1297 ), .b(
        \prgm_register/n1298 ), .out(\prgm_register/or_signal [648]) );
  nand2 \prgm_register/C5029  ( .a(enable), .b(a[648]), .out(
        \prgm_register/n1299 ) );
  nand2 \prgm_register/C5030  ( .a(\prgm_register/en_not ), .b(a[649]), .out(
        \prgm_register/n1300 ) );
  nand2 \prgm_register/C5031  ( .a(\prgm_register/n1299 ), .b(
        \prgm_register/n1300 ), .out(\prgm_register/or_signal [649]) );
  nand2 \prgm_register/C5032  ( .a(enable), .b(a[649]), .out(
        \prgm_register/n1301 ) );
  nand2 \prgm_register/C5033  ( .a(\prgm_register/en_not ), .b(a[650]), .out(
        \prgm_register/n1302 ) );
  nand2 \prgm_register/C5034  ( .a(\prgm_register/n1301 ), .b(
        \prgm_register/n1302 ), .out(\prgm_register/or_signal [650]) );
  nand2 \prgm_register/C5035  ( .a(enable), .b(a[650]), .out(
        \prgm_register/n1303 ) );
  nand2 \prgm_register/C5036  ( .a(\prgm_register/en_not ), .b(a[651]), .out(
        \prgm_register/n1304 ) );
  nand2 \prgm_register/C5037  ( .a(\prgm_register/n1303 ), .b(
        \prgm_register/n1304 ), .out(\prgm_register/or_signal [651]) );
  nand2 \prgm_register/C5038  ( .a(enable), .b(a[651]), .out(
        \prgm_register/n1305 ) );
  nand2 \prgm_register/C5039  ( .a(\prgm_register/en_not ), .b(a[652]), .out(
        \prgm_register/n1306 ) );
  nand2 \prgm_register/C5040  ( .a(\prgm_register/n1305 ), .b(
        \prgm_register/n1306 ), .out(\prgm_register/or_signal [652]) );
  nand2 \prgm_register/C5041  ( .a(enable), .b(a[652]), .out(
        \prgm_register/n1307 ) );
  nand2 \prgm_register/C5042  ( .a(\prgm_register/en_not ), .b(a[653]), .out(
        \prgm_register/n1308 ) );
  nand2 \prgm_register/C5043  ( .a(\prgm_register/n1307 ), .b(
        \prgm_register/n1308 ), .out(\prgm_register/or_signal [653]) );
  nand2 \prgm_register/C5044  ( .a(enable), .b(a[653]), .out(
        \prgm_register/n1309 ) );
  nand2 \prgm_register/C5045  ( .a(\prgm_register/en_not ), .b(a[654]), .out(
        \prgm_register/n1310 ) );
  nand2 \prgm_register/C5046  ( .a(\prgm_register/n1309 ), .b(
        \prgm_register/n1310 ), .out(\prgm_register/or_signal [654]) );
  nand2 \prgm_register/C5047  ( .a(enable), .b(a[654]), .out(
        \prgm_register/n1311 ) );
  nand2 \prgm_register/C5048  ( .a(\prgm_register/en_not ), .b(a[655]), .out(
        \prgm_register/n1312 ) );
  nand2 \prgm_register/C5049  ( .a(\prgm_register/n1311 ), .b(
        \prgm_register/n1312 ), .out(\prgm_register/or_signal [655]) );
  nand2 \prgm_register/C5050  ( .a(enable), .b(a[655]), .out(
        \prgm_register/n1313 ) );
  nand2 \prgm_register/C5051  ( .a(\prgm_register/en_not ), .b(a[656]), .out(
        \prgm_register/n1314 ) );
  nand2 \prgm_register/C5052  ( .a(\prgm_register/n1313 ), .b(
        \prgm_register/n1314 ), .out(\prgm_register/or_signal [656]) );
  nand2 \prgm_register/C5053  ( .a(enable), .b(a[656]), .out(
        \prgm_register/n1315 ) );
  nand2 \prgm_register/C5054  ( .a(\prgm_register/en_not ), .b(a[657]), .out(
        \prgm_register/n1316 ) );
  nand2 \prgm_register/C5055  ( .a(\prgm_register/n1315 ), .b(
        \prgm_register/n1316 ), .out(\prgm_register/or_signal [657]) );
  nand2 \prgm_register/C5056  ( .a(enable), .b(a[657]), .out(
        \prgm_register/n1317 ) );
  nand2 \prgm_register/C5057  ( .a(\prgm_register/en_not ), .b(a[658]), .out(
        \prgm_register/n1318 ) );
  nand2 \prgm_register/C5058  ( .a(\prgm_register/n1317 ), .b(
        \prgm_register/n1318 ), .out(\prgm_register/or_signal [658]) );
  nand2 \prgm_register/C5059  ( .a(enable), .b(a[658]), .out(
        \prgm_register/n1319 ) );
  nand2 \prgm_register/C5060  ( .a(\prgm_register/en_not ), .b(a[659]), .out(
        \prgm_register/n1320 ) );
  nand2 \prgm_register/C5061  ( .a(\prgm_register/n1319 ), .b(
        \prgm_register/n1320 ), .out(\prgm_register/or_signal [659]) );
  nand2 \prgm_register/C5062  ( .a(enable), .b(a[659]), .out(
        \prgm_register/n1321 ) );
  nand2 \prgm_register/C5063  ( .a(\prgm_register/en_not ), .b(a[660]), .out(
        \prgm_register/n1322 ) );
  nand2 \prgm_register/C5064  ( .a(\prgm_register/n1321 ), .b(
        \prgm_register/n1322 ), .out(\prgm_register/or_signal [660]) );
  nand2 \prgm_register/C5065  ( .a(enable), .b(a[660]), .out(
        \prgm_register/n1323 ) );
  nand2 \prgm_register/C5066  ( .a(\prgm_register/en_not ), .b(a[661]), .out(
        \prgm_register/n1324 ) );
  nand2 \prgm_register/C5067  ( .a(\prgm_register/n1323 ), .b(
        \prgm_register/n1324 ), .out(\prgm_register/or_signal [661]) );
  nand2 \prgm_register/C5068  ( .a(enable), .b(a[661]), .out(
        \prgm_register/n1325 ) );
  nand2 \prgm_register/C5069  ( .a(\prgm_register/en_not ), .b(a[662]), .out(
        \prgm_register/n1326 ) );
  nand2 \prgm_register/C5070  ( .a(\prgm_register/n1325 ), .b(
        \prgm_register/n1326 ), .out(\prgm_register/or_signal [662]) );
  nand2 \prgm_register/C5071  ( .a(enable), .b(a[662]), .out(
        \prgm_register/n1327 ) );
  nand2 \prgm_register/C5072  ( .a(\prgm_register/en_not ), .b(a[663]), .out(
        \prgm_register/n1328 ) );
  nand2 \prgm_register/C5073  ( .a(\prgm_register/n1327 ), .b(
        \prgm_register/n1328 ), .out(\prgm_register/or_signal [663]) );
  nand2 \prgm_register/C5074  ( .a(enable), .b(a[663]), .out(
        \prgm_register/n1329 ) );
  nand2 \prgm_register/C5075  ( .a(\prgm_register/en_not ), .b(a[664]), .out(
        \prgm_register/n1330 ) );
  nand2 \prgm_register/C5076  ( .a(\prgm_register/n1329 ), .b(
        \prgm_register/n1330 ), .out(\prgm_register/or_signal [664]) );
  nand2 \prgm_register/C5077  ( .a(enable), .b(a[664]), .out(
        \prgm_register/n1331 ) );
  nand2 \prgm_register/C5078  ( .a(\prgm_register/en_not ), .b(a[665]), .out(
        \prgm_register/n1332 ) );
  nand2 \prgm_register/C5079  ( .a(\prgm_register/n1331 ), .b(
        \prgm_register/n1332 ), .out(\prgm_register/or_signal [665]) );
  nand2 \prgm_register/C5080  ( .a(enable), .b(a[665]), .out(
        \prgm_register/n1333 ) );
  nand2 \prgm_register/C5081  ( .a(\prgm_register/en_not ), .b(a[666]), .out(
        \prgm_register/n1334 ) );
  nand2 \prgm_register/C5082  ( .a(\prgm_register/n1333 ), .b(
        \prgm_register/n1334 ), .out(\prgm_register/or_signal [666]) );
  nand2 \prgm_register/C5083  ( .a(enable), .b(a[666]), .out(
        \prgm_register/n1335 ) );
  nand2 \prgm_register/C5084  ( .a(\prgm_register/en_not ), .b(a[667]), .out(
        \prgm_register/n1336 ) );
  nand2 \prgm_register/C5085  ( .a(\prgm_register/n1335 ), .b(
        \prgm_register/n1336 ), .out(\prgm_register/or_signal [667]) );
  nand2 \prgm_register/C5086  ( .a(enable), .b(a[667]), .out(
        \prgm_register/n1337 ) );
  nand2 \prgm_register/C5087  ( .a(\prgm_register/en_not ), .b(a[668]), .out(
        \prgm_register/n1338 ) );
  nand2 \prgm_register/C5088  ( .a(\prgm_register/n1337 ), .b(
        \prgm_register/n1338 ), .out(\prgm_register/or_signal [668]) );
  nand2 \prgm_register/C5089  ( .a(enable), .b(a[668]), .out(
        \prgm_register/n1339 ) );
  nand2 \prgm_register/C5090  ( .a(\prgm_register/en_not ), .b(a[669]), .out(
        \prgm_register/n1340 ) );
  nand2 \prgm_register/C5091  ( .a(\prgm_register/n1339 ), .b(
        \prgm_register/n1340 ), .out(\prgm_register/or_signal [669]) );
  nand2 \prgm_register/C5092  ( .a(enable), .b(a[669]), .out(
        \prgm_register/n1341 ) );
  nand2 \prgm_register/C5093  ( .a(\prgm_register/en_not ), .b(a[670]), .out(
        \prgm_register/n1342 ) );
  nand2 \prgm_register/C5094  ( .a(\prgm_register/n1341 ), .b(
        \prgm_register/n1342 ), .out(\prgm_register/or_signal [670]) );
  nand2 \prgm_register/C5095  ( .a(enable), .b(a[670]), .out(
        \prgm_register/n1343 ) );
  nand2 \prgm_register/C5096  ( .a(\prgm_register/en_not ), .b(a[671]), .out(
        \prgm_register/n1344 ) );
  nand2 \prgm_register/C5097  ( .a(\prgm_register/n1343 ), .b(
        \prgm_register/n1344 ), .out(\prgm_register/or_signal [671]) );
  nand2 \prgm_register/C5098  ( .a(enable), .b(a[671]), .out(
        \prgm_register/n1345 ) );
  nand2 \prgm_register/C5099  ( .a(\prgm_register/en_not ), .b(a[672]), .out(
        \prgm_register/n1346 ) );
  nand2 \prgm_register/C5100  ( .a(\prgm_register/n1345 ), .b(
        \prgm_register/n1346 ), .out(\prgm_register/or_signal [672]) );
  nand2 \prgm_register/C5101  ( .a(enable), .b(a[672]), .out(
        \prgm_register/n1347 ) );
  nand2 \prgm_register/C5102  ( .a(\prgm_register/en_not ), .b(a[673]), .out(
        \prgm_register/n1348 ) );
  nand2 \prgm_register/C5103  ( .a(\prgm_register/n1347 ), .b(
        \prgm_register/n1348 ), .out(\prgm_register/or_signal [673]) );
  nand2 \prgm_register/C5104  ( .a(enable), .b(a[673]), .out(
        \prgm_register/n1349 ) );
  nand2 \prgm_register/C5105  ( .a(\prgm_register/en_not ), .b(a[674]), .out(
        \prgm_register/n1350 ) );
  nand2 \prgm_register/C5106  ( .a(\prgm_register/n1349 ), .b(
        \prgm_register/n1350 ), .out(\prgm_register/or_signal [674]) );
  nand2 \prgm_register/C5107  ( .a(enable), .b(a[674]), .out(
        \prgm_register/n1351 ) );
  nand2 \prgm_register/C5108  ( .a(\prgm_register/en_not ), .b(a[675]), .out(
        \prgm_register/n1352 ) );
  nand2 \prgm_register/C5109  ( .a(\prgm_register/n1351 ), .b(
        \prgm_register/n1352 ), .out(\prgm_register/or_signal [675]) );
  nand2 \prgm_register/C5110  ( .a(enable), .b(a[675]), .out(
        \prgm_register/n1353 ) );
  nand2 \prgm_register/C5111  ( .a(\prgm_register/en_not ), .b(a[676]), .out(
        \prgm_register/n1354 ) );
  nand2 \prgm_register/C5112  ( .a(\prgm_register/n1353 ), .b(
        \prgm_register/n1354 ), .out(\prgm_register/or_signal [676]) );
  nand2 \prgm_register/C5113  ( .a(enable), .b(a[676]), .out(
        \prgm_register/n1355 ) );
  nand2 \prgm_register/C5114  ( .a(\prgm_register/en_not ), .b(a[677]), .out(
        \prgm_register/n1356 ) );
  nand2 \prgm_register/C5115  ( .a(\prgm_register/n1355 ), .b(
        \prgm_register/n1356 ), .out(\prgm_register/or_signal [677]) );
  nand2 \prgm_register/C5116  ( .a(enable), .b(a[677]), .out(
        \prgm_register/n1357 ) );
  nand2 \prgm_register/C5117  ( .a(\prgm_register/en_not ), .b(a[678]), .out(
        \prgm_register/n1358 ) );
  nand2 \prgm_register/C5118  ( .a(\prgm_register/n1357 ), .b(
        \prgm_register/n1358 ), .out(\prgm_register/or_signal [678]) );
  nand2 \prgm_register/C5119  ( .a(enable), .b(a[678]), .out(
        \prgm_register/n1359 ) );
  nand2 \prgm_register/C5120  ( .a(\prgm_register/en_not ), .b(a[679]), .out(
        \prgm_register/n1360 ) );
  nand2 \prgm_register/C5121  ( .a(\prgm_register/n1359 ), .b(
        \prgm_register/n1360 ), .out(\prgm_register/or_signal [679]) );
  nand2 \prgm_register/C5122  ( .a(enable), .b(a[679]), .out(
        \prgm_register/n1361 ) );
  nand2 \prgm_register/C5123  ( .a(\prgm_register/en_not ), .b(a[680]), .out(
        \prgm_register/n1362 ) );
  nand2 \prgm_register/C5124  ( .a(\prgm_register/n1361 ), .b(
        \prgm_register/n1362 ), .out(\prgm_register/or_signal [680]) );
  nand2 \prgm_register/C5125  ( .a(enable), .b(a[680]), .out(
        \prgm_register/n1363 ) );
  nand2 \prgm_register/C5126  ( .a(\prgm_register/en_not ), .b(a[681]), .out(
        \prgm_register/n1364 ) );
  nand2 \prgm_register/C5127  ( .a(\prgm_register/n1363 ), .b(
        \prgm_register/n1364 ), .out(\prgm_register/or_signal [681]) );
  nand2 \prgm_register/C5128  ( .a(enable), .b(a[681]), .out(
        \prgm_register/n1365 ) );
  nand2 \prgm_register/C5129  ( .a(\prgm_register/en_not ), .b(a[682]), .out(
        \prgm_register/n1366 ) );
  nand2 \prgm_register/C5130  ( .a(\prgm_register/n1365 ), .b(
        \prgm_register/n1366 ), .out(\prgm_register/or_signal [682]) );
  nand2 \prgm_register/C5131  ( .a(enable), .b(a[682]), .out(
        \prgm_register/n1367 ) );
  nand2 \prgm_register/C5132  ( .a(\prgm_register/en_not ), .b(a[683]), .out(
        \prgm_register/n1368 ) );
  nand2 \prgm_register/C5133  ( .a(\prgm_register/n1367 ), .b(
        \prgm_register/n1368 ), .out(\prgm_register/or_signal [683]) );
  nand2 \prgm_register/C5134  ( .a(enable), .b(a[683]), .out(
        \prgm_register/n1369 ) );
  nand2 \prgm_register/C5135  ( .a(\prgm_register/en_not ), .b(a[684]), .out(
        \prgm_register/n1370 ) );
  nand2 \prgm_register/C5136  ( .a(\prgm_register/n1369 ), .b(
        \prgm_register/n1370 ), .out(\prgm_register/or_signal [684]) );
  nand2 \prgm_register/C5137  ( .a(enable), .b(a[684]), .out(
        \prgm_register/n1371 ) );
  nand2 \prgm_register/C5138  ( .a(\prgm_register/en_not ), .b(a[685]), .out(
        \prgm_register/n1372 ) );
  nand2 \prgm_register/C5139  ( .a(\prgm_register/n1371 ), .b(
        \prgm_register/n1372 ), .out(\prgm_register/or_signal [685]) );
  nand2 \prgm_register/C5140  ( .a(enable), .b(a[685]), .out(
        \prgm_register/n1373 ) );
  nand2 \prgm_register/C5141  ( .a(\prgm_register/en_not ), .b(a[686]), .out(
        \prgm_register/n1374 ) );
  nand2 \prgm_register/C5142  ( .a(\prgm_register/n1373 ), .b(
        \prgm_register/n1374 ), .out(\prgm_register/or_signal [686]) );
  nand2 \prgm_register/C5143  ( .a(enable), .b(a[686]), .out(
        \prgm_register/n1375 ) );
  nand2 \prgm_register/C5144  ( .a(\prgm_register/en_not ), .b(a[687]), .out(
        \prgm_register/n1376 ) );
  nand2 \prgm_register/C5145  ( .a(\prgm_register/n1375 ), .b(
        \prgm_register/n1376 ), .out(\prgm_register/or_signal [687]) );
  nand2 \prgm_register/C5146  ( .a(enable), .b(a[687]), .out(
        \prgm_register/n1377 ) );
  nand2 \prgm_register/C5147  ( .a(\prgm_register/en_not ), .b(a[688]), .out(
        \prgm_register/n1378 ) );
  nand2 \prgm_register/C5148  ( .a(\prgm_register/n1377 ), .b(
        \prgm_register/n1378 ), .out(\prgm_register/or_signal [688]) );
  nand2 \prgm_register/C5149  ( .a(enable), .b(a[688]), .out(
        \prgm_register/n1379 ) );
  nand2 \prgm_register/C5150  ( .a(\prgm_register/en_not ), .b(a[689]), .out(
        \prgm_register/n1380 ) );
  nand2 \prgm_register/C5151  ( .a(\prgm_register/n1379 ), .b(
        \prgm_register/n1380 ), .out(\prgm_register/or_signal [689]) );
  nand2 \prgm_register/C5152  ( .a(enable), .b(a[689]), .out(
        \prgm_register/n1381 ) );
  nand2 \prgm_register/C5153  ( .a(\prgm_register/en_not ), .b(a[690]), .out(
        \prgm_register/n1382 ) );
  nand2 \prgm_register/C5154  ( .a(\prgm_register/n1381 ), .b(
        \prgm_register/n1382 ), .out(\prgm_register/or_signal [690]) );
  nand2 \prgm_register/C5155  ( .a(enable), .b(a[690]), .out(
        \prgm_register/n1383 ) );
  nand2 \prgm_register/C5156  ( .a(\prgm_register/en_not ), .b(a[691]), .out(
        \prgm_register/n1384 ) );
  nand2 \prgm_register/C5157  ( .a(\prgm_register/n1383 ), .b(
        \prgm_register/n1384 ), .out(\prgm_register/or_signal [691]) );
  nand2 \prgm_register/C5158  ( .a(enable), .b(a[691]), .out(
        \prgm_register/n1385 ) );
  nand2 \prgm_register/C5159  ( .a(\prgm_register/en_not ), .b(a[692]), .out(
        \prgm_register/n1386 ) );
  nand2 \prgm_register/C5160  ( .a(\prgm_register/n1385 ), .b(
        \prgm_register/n1386 ), .out(\prgm_register/or_signal [692]) );
  nand2 \prgm_register/C5161  ( .a(enable), .b(a[692]), .out(
        \prgm_register/n1387 ) );
  nand2 \prgm_register/C5162  ( .a(\prgm_register/en_not ), .b(a[693]), .out(
        \prgm_register/n1388 ) );
  nand2 \prgm_register/C5163  ( .a(\prgm_register/n1387 ), .b(
        \prgm_register/n1388 ), .out(\prgm_register/or_signal [693]) );
  nand2 \prgm_register/C5164  ( .a(enable), .b(a[693]), .out(
        \prgm_register/n1389 ) );
  nand2 \prgm_register/C5165  ( .a(\prgm_register/en_not ), .b(a[694]), .out(
        \prgm_register/n1390 ) );
  nand2 \prgm_register/C5166  ( .a(\prgm_register/n1389 ), .b(
        \prgm_register/n1390 ), .out(\prgm_register/or_signal [694]) );
  nand2 \prgm_register/C5167  ( .a(enable), .b(a[694]), .out(
        \prgm_register/n1391 ) );
  nand2 \prgm_register/C5168  ( .a(\prgm_register/en_not ), .b(a[695]), .out(
        \prgm_register/n1392 ) );
  nand2 \prgm_register/C5169  ( .a(\prgm_register/n1391 ), .b(
        \prgm_register/n1392 ), .out(\prgm_register/or_signal [695]) );
  nand2 \prgm_register/C5170  ( .a(enable), .b(a[695]), .out(
        \prgm_register/n1393 ) );
  nand2 \prgm_register/C5171  ( .a(\prgm_register/en_not ), .b(a[696]), .out(
        \prgm_register/n1394 ) );
  nand2 \prgm_register/C5172  ( .a(\prgm_register/n1393 ), .b(
        \prgm_register/n1394 ), .out(\prgm_register/or_signal [696]) );
  nand2 \prgm_register/C5173  ( .a(enable), .b(a[696]), .out(
        \prgm_register/n1395 ) );
  nand2 \prgm_register/C5174  ( .a(\prgm_register/en_not ), .b(a[697]), .out(
        \prgm_register/n1396 ) );
  nand2 \prgm_register/C5175  ( .a(\prgm_register/n1395 ), .b(
        \prgm_register/n1396 ), .out(\prgm_register/or_signal [697]) );
  nand2 \prgm_register/C5176  ( .a(enable), .b(a[697]), .out(
        \prgm_register/n1397 ) );
  nand2 \prgm_register/C5177  ( .a(\prgm_register/en_not ), .b(a[698]), .out(
        \prgm_register/n1398 ) );
  nand2 \prgm_register/C5178  ( .a(\prgm_register/n1397 ), .b(
        \prgm_register/n1398 ), .out(\prgm_register/or_signal [698]) );
  nand2 \prgm_register/C5179  ( .a(enable), .b(a[698]), .out(
        \prgm_register/n1399 ) );
  nand2 \prgm_register/C5180  ( .a(\prgm_register/en_not ), .b(a[699]), .out(
        \prgm_register/n1400 ) );
  nand2 \prgm_register/C5181  ( .a(\prgm_register/n1399 ), .b(
        \prgm_register/n1400 ), .out(\prgm_register/or_signal [699]) );
  nand2 \prgm_register/C5182  ( .a(enable), .b(a[699]), .out(
        \prgm_register/n1401 ) );
  nand2 \prgm_register/C5183  ( .a(\prgm_register/en_not ), .b(a[700]), .out(
        \prgm_register/n1402 ) );
  nand2 \prgm_register/C5184  ( .a(\prgm_register/n1401 ), .b(
        \prgm_register/n1402 ), .out(\prgm_register/or_signal [700]) );
  nand2 \prgm_register/C5185  ( .a(enable), .b(a[700]), .out(
        \prgm_register/n1403 ) );
  nand2 \prgm_register/C5186  ( .a(\prgm_register/en_not ), .b(a[701]), .out(
        \prgm_register/n1404 ) );
  nand2 \prgm_register/C5187  ( .a(\prgm_register/n1403 ), .b(
        \prgm_register/n1404 ), .out(\prgm_register/or_signal [701]) );
  nand2 \prgm_register/C5188  ( .a(enable), .b(a[701]), .out(
        \prgm_register/n1405 ) );
  nand2 \prgm_register/C5189  ( .a(\prgm_register/en_not ), .b(a[702]), .out(
        \prgm_register/n1406 ) );
  nand2 \prgm_register/C5190  ( .a(\prgm_register/n1405 ), .b(
        \prgm_register/n1406 ), .out(\prgm_register/or_signal [702]) );
  nand2 \prgm_register/C5191  ( .a(enable), .b(a[702]), .out(
        \prgm_register/n1407 ) );
  nand2 \prgm_register/C5192  ( .a(\prgm_register/en_not ), .b(a[703]), .out(
        \prgm_register/n1408 ) );
  nand2 \prgm_register/C5193  ( .a(\prgm_register/n1407 ), .b(
        \prgm_register/n1408 ), .out(\prgm_register/or_signal [703]) );
  nand2 \prgm_register/C5194  ( .a(enable), .b(a[703]), .out(
        \prgm_register/n1409 ) );
  nand2 \prgm_register/C5195  ( .a(\prgm_register/en_not ), .b(a[704]), .out(
        \prgm_register/n1410 ) );
  nand2 \prgm_register/C5196  ( .a(\prgm_register/n1409 ), .b(
        \prgm_register/n1410 ), .out(\prgm_register/or_signal [704]) );
  nand2 \prgm_register/C5197  ( .a(enable), .b(a[704]), .out(
        \prgm_register/n1411 ) );
  nand2 \prgm_register/C5198  ( .a(\prgm_register/en_not ), .b(a[705]), .out(
        \prgm_register/n1412 ) );
  nand2 \prgm_register/C5199  ( .a(\prgm_register/n1411 ), .b(
        \prgm_register/n1412 ), .out(\prgm_register/or_signal [705]) );
  nand2 \prgm_register/C5200  ( .a(enable), .b(a[705]), .out(
        \prgm_register/n1413 ) );
  nand2 \prgm_register/C5201  ( .a(\prgm_register/en_not ), .b(a[706]), .out(
        \prgm_register/n1414 ) );
  nand2 \prgm_register/C5202  ( .a(\prgm_register/n1413 ), .b(
        \prgm_register/n1414 ), .out(\prgm_register/or_signal [706]) );
  nand2 \prgm_register/C5203  ( .a(enable), .b(a[706]), .out(
        \prgm_register/n1415 ) );
  nand2 \prgm_register/C5204  ( .a(\prgm_register/en_not ), .b(a[707]), .out(
        \prgm_register/n1416 ) );
  nand2 \prgm_register/C5205  ( .a(\prgm_register/n1415 ), .b(
        \prgm_register/n1416 ), .out(\prgm_register/or_signal [707]) );
  nand2 \prgm_register/C5206  ( .a(enable), .b(a[707]), .out(
        \prgm_register/n1417 ) );
  nand2 \prgm_register/C5207  ( .a(\prgm_register/en_not ), .b(a[708]), .out(
        \prgm_register/n1418 ) );
  nand2 \prgm_register/C5208  ( .a(\prgm_register/n1417 ), .b(
        \prgm_register/n1418 ), .out(\prgm_register/or_signal [708]) );
  nand2 \prgm_register/C5209  ( .a(enable), .b(a[708]), .out(
        \prgm_register/n1419 ) );
  nand2 \prgm_register/C5210  ( .a(\prgm_register/en_not ), .b(a[709]), .out(
        \prgm_register/n1420 ) );
  nand2 \prgm_register/C5211  ( .a(\prgm_register/n1419 ), .b(
        \prgm_register/n1420 ), .out(\prgm_register/or_signal [709]) );
  nand2 \prgm_register/C5212  ( .a(enable), .b(a[709]), .out(
        \prgm_register/n1421 ) );
  nand2 \prgm_register/C5213  ( .a(\prgm_register/en_not ), .b(a[710]), .out(
        \prgm_register/n1422 ) );
  nand2 \prgm_register/C5214  ( .a(\prgm_register/n1421 ), .b(
        \prgm_register/n1422 ), .out(\prgm_register/or_signal [710]) );
  nand2 \prgm_register/C5215  ( .a(enable), .b(a[710]), .out(
        \prgm_register/n1423 ) );
  nand2 \prgm_register/C5216  ( .a(\prgm_register/en_not ), .b(a[711]), .out(
        \prgm_register/n1424 ) );
  nand2 \prgm_register/C5217  ( .a(\prgm_register/n1423 ), .b(
        \prgm_register/n1424 ), .out(\prgm_register/or_signal [711]) );
  nand2 \prgm_register/C5218  ( .a(enable), .b(a[711]), .out(
        \prgm_register/n1425 ) );
  nand2 \prgm_register/C5219  ( .a(\prgm_register/en_not ), .b(a[712]), .out(
        \prgm_register/n1426 ) );
  nand2 \prgm_register/C5220  ( .a(\prgm_register/n1425 ), .b(
        \prgm_register/n1426 ), .out(\prgm_register/or_signal [712]) );
  nand2 \prgm_register/C5221  ( .a(enable), .b(a[712]), .out(
        \prgm_register/n1427 ) );
  nand2 \prgm_register/C5222  ( .a(\prgm_register/en_not ), .b(a[713]), .out(
        \prgm_register/n1428 ) );
  nand2 \prgm_register/C5223  ( .a(\prgm_register/n1427 ), .b(
        \prgm_register/n1428 ), .out(\prgm_register/or_signal [713]) );
  nand2 \prgm_register/C5224  ( .a(enable), .b(a[713]), .out(
        \prgm_register/n1429 ) );
  nand2 \prgm_register/C5225  ( .a(\prgm_register/en_not ), .b(a[714]), .out(
        \prgm_register/n1430 ) );
  nand2 \prgm_register/C5226  ( .a(\prgm_register/n1429 ), .b(
        \prgm_register/n1430 ), .out(\prgm_register/or_signal [714]) );
  nand2 \prgm_register/C5227  ( .a(enable), .b(a[714]), .out(
        \prgm_register/n1431 ) );
  nand2 \prgm_register/C5228  ( .a(\prgm_register/en_not ), .b(a[715]), .out(
        \prgm_register/n1432 ) );
  nand2 \prgm_register/C5229  ( .a(\prgm_register/n1431 ), .b(
        \prgm_register/n1432 ), .out(\prgm_register/or_signal [715]) );
  nand2 \prgm_register/C5230  ( .a(enable), .b(a[715]), .out(
        \prgm_register/n1433 ) );
  nand2 \prgm_register/C5231  ( .a(\prgm_register/en_not ), .b(a[716]), .out(
        \prgm_register/n1434 ) );
  nand2 \prgm_register/C5232  ( .a(\prgm_register/n1433 ), .b(
        \prgm_register/n1434 ), .out(\prgm_register/or_signal [716]) );
  nand2 \prgm_register/C5233  ( .a(enable), .b(a[716]), .out(
        \prgm_register/n1435 ) );
  nand2 \prgm_register/C5234  ( .a(\prgm_register/en_not ), .b(a[717]), .out(
        \prgm_register/n1436 ) );
  nand2 \prgm_register/C5235  ( .a(\prgm_register/n1435 ), .b(
        \prgm_register/n1436 ), .out(\prgm_register/or_signal [717]) );
  nand2 \prgm_register/C5236  ( .a(enable), .b(a[717]), .out(
        \prgm_register/n1437 ) );
  nand2 \prgm_register/C5237  ( .a(\prgm_register/en_not ), .b(a[718]), .out(
        \prgm_register/n1438 ) );
  nand2 \prgm_register/C5238  ( .a(\prgm_register/n1437 ), .b(
        \prgm_register/n1438 ), .out(\prgm_register/or_signal [718]) );
  nand2 \prgm_register/C5239  ( .a(enable), .b(a[718]), .out(
        \prgm_register/n1439 ) );
  nand2 \prgm_register/C5240  ( .a(\prgm_register/en_not ), .b(a[719]), .out(
        \prgm_register/n1440 ) );
  nand2 \prgm_register/C5241  ( .a(\prgm_register/n1439 ), .b(
        \prgm_register/n1440 ), .out(\prgm_register/or_signal [719]) );
  nand2 \prgm_register/C5242  ( .a(enable), .b(a[719]), .out(
        \prgm_register/n1441 ) );
  nand2 \prgm_register/C5243  ( .a(\prgm_register/en_not ), .b(a[720]), .out(
        \prgm_register/n1442 ) );
  nand2 \prgm_register/C5244  ( .a(\prgm_register/n1441 ), .b(
        \prgm_register/n1442 ), .out(\prgm_register/or_signal [720]) );
  nand2 \prgm_register/C5245  ( .a(enable), .b(a[720]), .out(
        \prgm_register/n1443 ) );
  nand2 \prgm_register/C5246  ( .a(\prgm_register/en_not ), .b(a[721]), .out(
        \prgm_register/n1444 ) );
  nand2 \prgm_register/C5247  ( .a(\prgm_register/n1443 ), .b(
        \prgm_register/n1444 ), .out(\prgm_register/or_signal [721]) );
  nand2 \prgm_register/C5248  ( .a(enable), .b(a[721]), .out(
        \prgm_register/n1445 ) );
  nand2 \prgm_register/C5249  ( .a(\prgm_register/en_not ), .b(a[722]), .out(
        \prgm_register/n1446 ) );
  nand2 \prgm_register/C5250  ( .a(\prgm_register/n1445 ), .b(
        \prgm_register/n1446 ), .out(\prgm_register/or_signal [722]) );
  nand2 \prgm_register/C5251  ( .a(enable), .b(a[722]), .out(
        \prgm_register/n1447 ) );
  nand2 \prgm_register/C5252  ( .a(\prgm_register/en_not ), .b(a[723]), .out(
        \prgm_register/n1448 ) );
  nand2 \prgm_register/C5253  ( .a(\prgm_register/n1447 ), .b(
        \prgm_register/n1448 ), .out(\prgm_register/or_signal [723]) );
  nand2 \prgm_register/C5254  ( .a(enable), .b(a[723]), .out(
        \prgm_register/n1449 ) );
  nand2 \prgm_register/C5255  ( .a(\prgm_register/en_not ), .b(a[724]), .out(
        \prgm_register/n1450 ) );
  nand2 \prgm_register/C5256  ( .a(\prgm_register/n1449 ), .b(
        \prgm_register/n1450 ), .out(\prgm_register/or_signal [724]) );
  nand2 \prgm_register/C5257  ( .a(enable), .b(a[724]), .out(
        \prgm_register/n1451 ) );
  nand2 \prgm_register/C5258  ( .a(\prgm_register/en_not ), .b(a[725]), .out(
        \prgm_register/n1452 ) );
  nand2 \prgm_register/C5259  ( .a(\prgm_register/n1451 ), .b(
        \prgm_register/n1452 ), .out(\prgm_register/or_signal [725]) );
  nand2 \prgm_register/C5260  ( .a(enable), .b(a[725]), .out(
        \prgm_register/n1453 ) );
  nand2 \prgm_register/C5261  ( .a(\prgm_register/en_not ), .b(a[726]), .out(
        \prgm_register/n1454 ) );
  nand2 \prgm_register/C5262  ( .a(\prgm_register/n1453 ), .b(
        \prgm_register/n1454 ), .out(\prgm_register/or_signal [726]) );
  nand2 \prgm_register/C5263  ( .a(enable), .b(a[726]), .out(
        \prgm_register/n1455 ) );
  nand2 \prgm_register/C5264  ( .a(\prgm_register/en_not ), .b(a[727]), .out(
        \prgm_register/n1456 ) );
  nand2 \prgm_register/C5265  ( .a(\prgm_register/n1455 ), .b(
        \prgm_register/n1456 ), .out(\prgm_register/or_signal [727]) );
  nand2 \prgm_register/C5266  ( .a(enable), .b(a[727]), .out(
        \prgm_register/n1457 ) );
  nand2 \prgm_register/C5267  ( .a(\prgm_register/en_not ), .b(a[728]), .out(
        \prgm_register/n1458 ) );
  nand2 \prgm_register/C5268  ( .a(\prgm_register/n1457 ), .b(
        \prgm_register/n1458 ), .out(\prgm_register/or_signal [728]) );
  nand2 \prgm_register/C5269  ( .a(enable), .b(a[728]), .out(
        \prgm_register/n1459 ) );
  nand2 \prgm_register/C5270  ( .a(\prgm_register/en_not ), .b(a[729]), .out(
        \prgm_register/n1460 ) );
  nand2 \prgm_register/C5271  ( .a(\prgm_register/n1459 ), .b(
        \prgm_register/n1460 ), .out(\prgm_register/or_signal [729]) );
  nand2 \prgm_register/C5272  ( .a(enable), .b(a[729]), .out(
        \prgm_register/n1461 ) );
  nand2 \prgm_register/C5273  ( .a(\prgm_register/en_not ), .b(a[730]), .out(
        \prgm_register/n1462 ) );
  nand2 \prgm_register/C5274  ( .a(\prgm_register/n1461 ), .b(
        \prgm_register/n1462 ), .out(\prgm_register/or_signal [730]) );
  nand2 \prgm_register/C5275  ( .a(enable), .b(a[730]), .out(
        \prgm_register/n1463 ) );
  nand2 \prgm_register/C5276  ( .a(\prgm_register/en_not ), .b(a[731]), .out(
        \prgm_register/n1464 ) );
  nand2 \prgm_register/C5277  ( .a(\prgm_register/n1463 ), .b(
        \prgm_register/n1464 ), .out(\prgm_register/or_signal [731]) );
  nand2 \prgm_register/C5278  ( .a(enable), .b(a[731]), .out(
        \prgm_register/n1465 ) );
  nand2 \prgm_register/C5279  ( .a(\prgm_register/en_not ), .b(a[732]), .out(
        \prgm_register/n1466 ) );
  nand2 \prgm_register/C5280  ( .a(\prgm_register/n1465 ), .b(
        \prgm_register/n1466 ), .out(\prgm_register/or_signal [732]) );
  nand2 \prgm_register/C5281  ( .a(enable), .b(a[732]), .out(
        \prgm_register/n1467 ) );
  nand2 \prgm_register/C5282  ( .a(\prgm_register/en_not ), .b(a[733]), .out(
        \prgm_register/n1468 ) );
  nand2 \prgm_register/C5283  ( .a(\prgm_register/n1467 ), .b(
        \prgm_register/n1468 ), .out(\prgm_register/or_signal [733]) );
  nand2 \prgm_register/C5284  ( .a(enable), .b(a[733]), .out(
        \prgm_register/n1469 ) );
  nand2 \prgm_register/C5285  ( .a(\prgm_register/en_not ), .b(a[734]), .out(
        \prgm_register/n1470 ) );
  nand2 \prgm_register/C5286  ( .a(\prgm_register/n1469 ), .b(
        \prgm_register/n1470 ), .out(\prgm_register/or_signal [734]) );
  nand2 \prgm_register/C5287  ( .a(enable), .b(a[734]), .out(
        \prgm_register/n1471 ) );
  nand2 \prgm_register/C5288  ( .a(\prgm_register/en_not ), .b(a[735]), .out(
        \prgm_register/n1472 ) );
  nand2 \prgm_register/C5289  ( .a(\prgm_register/n1471 ), .b(
        \prgm_register/n1472 ), .out(\prgm_register/or_signal [735]) );
  nand2 \prgm_register/C5290  ( .a(enable), .b(a[735]), .out(
        \prgm_register/n1473 ) );
  nand2 \prgm_register/C5291  ( .a(\prgm_register/en_not ), .b(a[736]), .out(
        \prgm_register/n1474 ) );
  nand2 \prgm_register/C5292  ( .a(\prgm_register/n1473 ), .b(
        \prgm_register/n1474 ), .out(\prgm_register/or_signal [736]) );
  nand2 \prgm_register/C5293  ( .a(enable), .b(a[736]), .out(
        \prgm_register/n1475 ) );
  nand2 \prgm_register/C5294  ( .a(\prgm_register/en_not ), .b(a[737]), .out(
        \prgm_register/n1476 ) );
  nand2 \prgm_register/C5295  ( .a(\prgm_register/n1475 ), .b(
        \prgm_register/n1476 ), .out(\prgm_register/or_signal [737]) );
  nand2 \prgm_register/C5296  ( .a(enable), .b(a[737]), .out(
        \prgm_register/n1477 ) );
  nand2 \prgm_register/C5297  ( .a(\prgm_register/en_not ), .b(a[738]), .out(
        \prgm_register/n1478 ) );
  nand2 \prgm_register/C5298  ( .a(\prgm_register/n1477 ), .b(
        \prgm_register/n1478 ), .out(\prgm_register/or_signal [738]) );
  nand2 \prgm_register/C5299  ( .a(enable), .b(a[738]), .out(
        \prgm_register/n1479 ) );
  nand2 \prgm_register/C5300  ( .a(\prgm_register/en_not ), .b(a[739]), .out(
        \prgm_register/n1480 ) );
  nand2 \prgm_register/C5301  ( .a(\prgm_register/n1479 ), .b(
        \prgm_register/n1480 ), .out(\prgm_register/or_signal [739]) );
  nand2 \prgm_register/C5302  ( .a(enable), .b(a[739]), .out(
        \prgm_register/n1481 ) );
  nand2 \prgm_register/C5303  ( .a(\prgm_register/en_not ), .b(a[740]), .out(
        \prgm_register/n1482 ) );
  nand2 \prgm_register/C5304  ( .a(\prgm_register/n1481 ), .b(
        \prgm_register/n1482 ), .out(\prgm_register/or_signal [740]) );
  nand2 \prgm_register/C5305  ( .a(enable), .b(a[740]), .out(
        \prgm_register/n1483 ) );
  nand2 \prgm_register/C5306  ( .a(\prgm_register/en_not ), .b(a[741]), .out(
        \prgm_register/n1484 ) );
  nand2 \prgm_register/C5307  ( .a(\prgm_register/n1483 ), .b(
        \prgm_register/n1484 ), .out(\prgm_register/or_signal [741]) );
  nand2 \prgm_register/C5308  ( .a(enable), .b(a[741]), .out(
        \prgm_register/n1485 ) );
  nand2 \prgm_register/C5309  ( .a(\prgm_register/en_not ), .b(a[742]), .out(
        \prgm_register/n1486 ) );
  nand2 \prgm_register/C5310  ( .a(\prgm_register/n1485 ), .b(
        \prgm_register/n1486 ), .out(\prgm_register/or_signal [742]) );
  nand2 \prgm_register/C5311  ( .a(enable), .b(a[742]), .out(
        \prgm_register/n1487 ) );
  nand2 \prgm_register/C5312  ( .a(\prgm_register/en_not ), .b(a[743]), .out(
        \prgm_register/n1488 ) );
  nand2 \prgm_register/C5313  ( .a(\prgm_register/n1487 ), .b(
        \prgm_register/n1488 ), .out(\prgm_register/or_signal [743]) );
  nand2 \prgm_register/C5314  ( .a(enable), .b(a[743]), .out(
        \prgm_register/n1489 ) );
  nand2 \prgm_register/C5315  ( .a(\prgm_register/en_not ), .b(a[744]), .out(
        \prgm_register/n1490 ) );
  nand2 \prgm_register/C5316  ( .a(\prgm_register/n1489 ), .b(
        \prgm_register/n1490 ), .out(\prgm_register/or_signal [744]) );
  nand2 \prgm_register/C5317  ( .a(enable), .b(a[744]), .out(
        \prgm_register/n1491 ) );
  nand2 \prgm_register/C5318  ( .a(\prgm_register/en_not ), .b(a[745]), .out(
        \prgm_register/n1492 ) );
  nand2 \prgm_register/C5319  ( .a(\prgm_register/n1491 ), .b(
        \prgm_register/n1492 ), .out(\prgm_register/or_signal [745]) );
  nand2 \prgm_register/C5320  ( .a(enable), .b(a[745]), .out(
        \prgm_register/n1493 ) );
  nand2 \prgm_register/C5321  ( .a(\prgm_register/en_not ), .b(a[746]), .out(
        \prgm_register/n1494 ) );
  nand2 \prgm_register/C5322  ( .a(\prgm_register/n1493 ), .b(
        \prgm_register/n1494 ), .out(\prgm_register/or_signal [746]) );
  nand2 \prgm_register/C5323  ( .a(enable), .b(a[746]), .out(
        \prgm_register/n1495 ) );
  nand2 \prgm_register/C5324  ( .a(\prgm_register/en_not ), .b(a[747]), .out(
        \prgm_register/n1496 ) );
  nand2 \prgm_register/C5325  ( .a(\prgm_register/n1495 ), .b(
        \prgm_register/n1496 ), .out(\prgm_register/or_signal [747]) );
  nand2 \prgm_register/C5326  ( .a(enable), .b(a[747]), .out(
        \prgm_register/n1497 ) );
  nand2 \prgm_register/C5327  ( .a(\prgm_register/en_not ), .b(a[748]), .out(
        \prgm_register/n1498 ) );
  nand2 \prgm_register/C5328  ( .a(\prgm_register/n1497 ), .b(
        \prgm_register/n1498 ), .out(\prgm_register/or_signal [748]) );
  nand2 \prgm_register/C5329  ( .a(enable), .b(a[748]), .out(
        \prgm_register/n1499 ) );
  nand2 \prgm_register/C5330  ( .a(\prgm_register/en_not ), .b(a[749]), .out(
        \prgm_register/n1500 ) );
  nand2 \prgm_register/C5331  ( .a(\prgm_register/n1499 ), .b(
        \prgm_register/n1500 ), .out(\prgm_register/or_signal [749]) );
  nand2 \prgm_register/C5332  ( .a(enable), .b(a[749]), .out(
        \prgm_register/n1501 ) );
  nand2 \prgm_register/C5333  ( .a(\prgm_register/en_not ), .b(a[750]), .out(
        \prgm_register/n1502 ) );
  nand2 \prgm_register/C5334  ( .a(\prgm_register/n1501 ), .b(
        \prgm_register/n1502 ), .out(\prgm_register/or_signal [750]) );
  nand2 \prgm_register/C5335  ( .a(enable), .b(a[750]), .out(
        \prgm_register/n1503 ) );
  nand2 \prgm_register/C5336  ( .a(\prgm_register/en_not ), .b(a[751]), .out(
        \prgm_register/n1504 ) );
  nand2 \prgm_register/C5337  ( .a(\prgm_register/n1503 ), .b(
        \prgm_register/n1504 ), .out(\prgm_register/or_signal [751]) );
  nand2 \prgm_register/C5338  ( .a(enable), .b(a[751]), .out(
        \prgm_register/n1505 ) );
  nand2 \prgm_register/C5339  ( .a(\prgm_register/en_not ), .b(a[752]), .out(
        \prgm_register/n1506 ) );
  nand2 \prgm_register/C5340  ( .a(\prgm_register/n1505 ), .b(
        \prgm_register/n1506 ), .out(\prgm_register/or_signal [752]) );
  nand2 \prgm_register/C5341  ( .a(enable), .b(a[752]), .out(
        \prgm_register/n1507 ) );
  nand2 \prgm_register/C5342  ( .a(\prgm_register/en_not ), .b(a[753]), .out(
        \prgm_register/n1508 ) );
  nand2 \prgm_register/C5343  ( .a(\prgm_register/n1507 ), .b(
        \prgm_register/n1508 ), .out(\prgm_register/or_signal [753]) );
  nand2 \prgm_register/C5344  ( .a(enable), .b(a[753]), .out(
        \prgm_register/n1509 ) );
  nand2 \prgm_register/C5345  ( .a(\prgm_register/en_not ), .b(a[754]), .out(
        \prgm_register/n1510 ) );
  nand2 \prgm_register/C5346  ( .a(\prgm_register/n1509 ), .b(
        \prgm_register/n1510 ), .out(\prgm_register/or_signal [754]) );
  nand2 \prgm_register/C5347  ( .a(enable), .b(a[754]), .out(
        \prgm_register/n1511 ) );
  nand2 \prgm_register/C5348  ( .a(\prgm_register/en_not ), .b(a[755]), .out(
        \prgm_register/n1512 ) );
  nand2 \prgm_register/C5349  ( .a(\prgm_register/n1511 ), .b(
        \prgm_register/n1512 ), .out(\prgm_register/or_signal [755]) );
  nand2 \prgm_register/C5350  ( .a(enable), .b(a[755]), .out(
        \prgm_register/n1513 ) );
  nand2 \prgm_register/C5351  ( .a(\prgm_register/en_not ), .b(a[756]), .out(
        \prgm_register/n1514 ) );
  nand2 \prgm_register/C5352  ( .a(\prgm_register/n1513 ), .b(
        \prgm_register/n1514 ), .out(\prgm_register/or_signal [756]) );
  nand2 \prgm_register/C5353  ( .a(enable), .b(a[756]), .out(
        \prgm_register/n1515 ) );
  nand2 \prgm_register/C5354  ( .a(\prgm_register/en_not ), .b(a[757]), .out(
        \prgm_register/n1516 ) );
  nand2 \prgm_register/C5355  ( .a(\prgm_register/n1515 ), .b(
        \prgm_register/n1516 ), .out(\prgm_register/or_signal [757]) );
  nand2 \prgm_register/C5356  ( .a(enable), .b(a[757]), .out(
        \prgm_register/n1517 ) );
  nand2 \prgm_register/C5357  ( .a(\prgm_register/en_not ), .b(a[758]), .out(
        \prgm_register/n1518 ) );
  nand2 \prgm_register/C5358  ( .a(\prgm_register/n1517 ), .b(
        \prgm_register/n1518 ), .out(\prgm_register/or_signal [758]) );
  nand2 \prgm_register/C5359  ( .a(enable), .b(a[758]), .out(
        \prgm_register/n1519 ) );
  nand2 \prgm_register/C5360  ( .a(\prgm_register/en_not ), .b(a[759]), .out(
        \prgm_register/n1520 ) );
  nand2 \prgm_register/C5361  ( .a(\prgm_register/n1519 ), .b(
        \prgm_register/n1520 ), .out(\prgm_register/or_signal [759]) );
  nand2 \prgm_register/C5362  ( .a(enable), .b(a[759]), .out(
        \prgm_register/n1521 ) );
  nand2 \prgm_register/C5363  ( .a(\prgm_register/en_not ), .b(a[760]), .out(
        \prgm_register/n1522 ) );
  nand2 \prgm_register/C5364  ( .a(\prgm_register/n1521 ), .b(
        \prgm_register/n1522 ), .out(\prgm_register/or_signal [760]) );
  nand2 \prgm_register/C5365  ( .a(enable), .b(a[760]), .out(
        \prgm_register/n1523 ) );
  nand2 \prgm_register/C5366  ( .a(\prgm_register/en_not ), .b(a[761]), .out(
        \prgm_register/n1524 ) );
  nand2 \prgm_register/C5367  ( .a(\prgm_register/n1523 ), .b(
        \prgm_register/n1524 ), .out(\prgm_register/or_signal [761]) );
  nand2 \prgm_register/C5368  ( .a(enable), .b(a[761]), .out(
        \prgm_register/n1525 ) );
  nand2 \prgm_register/C5369  ( .a(\prgm_register/en_not ), .b(a[762]), .out(
        \prgm_register/n1526 ) );
  nand2 \prgm_register/C5370  ( .a(\prgm_register/n1525 ), .b(
        \prgm_register/n1526 ), .out(\prgm_register/or_signal [762]) );
  nand2 \prgm_register/C5371  ( .a(enable), .b(a[762]), .out(
        \prgm_register/n1527 ) );
  nand2 \prgm_register/C5372  ( .a(\prgm_register/en_not ), .b(a[763]), .out(
        \prgm_register/n1528 ) );
  nand2 \prgm_register/C5373  ( .a(\prgm_register/n1527 ), .b(
        \prgm_register/n1528 ), .out(\prgm_register/or_signal [763]) );
  nand2 \prgm_register/C5374  ( .a(enable), .b(a[763]), .out(
        \prgm_register/n1529 ) );
  nand2 \prgm_register/C5375  ( .a(\prgm_register/en_not ), .b(a[764]), .out(
        \prgm_register/n1530 ) );
  nand2 \prgm_register/C5376  ( .a(\prgm_register/n1529 ), .b(
        \prgm_register/n1530 ), .out(\prgm_register/or_signal [764]) );
  nand2 \prgm_register/C5377  ( .a(enable), .b(a[764]), .out(
        \prgm_register/n1531 ) );
  nand2 \prgm_register/C5378  ( .a(\prgm_register/en_not ), .b(a[765]), .out(
        \prgm_register/n1532 ) );
  nand2 \prgm_register/C5379  ( .a(\prgm_register/n1531 ), .b(
        \prgm_register/n1532 ), .out(\prgm_register/or_signal [765]) );
  nand2 \prgm_register/C5380  ( .a(enable), .b(a[765]), .out(
        \prgm_register/n1533 ) );
  nand2 \prgm_register/C5381  ( .a(\prgm_register/en_not ), .b(a[766]), .out(
        \prgm_register/n1534 ) );
  nand2 \prgm_register/C5382  ( .a(\prgm_register/n1533 ), .b(
        \prgm_register/n1534 ), .out(\prgm_register/or_signal [766]) );
  nand2 \prgm_register/C5383  ( .a(enable), .b(a[766]), .out(
        \prgm_register/n1535 ) );
  nand2 \prgm_register/C5384  ( .a(\prgm_register/en_not ), .b(a[767]), .out(
        \prgm_register/n1536 ) );
  nand2 \prgm_register/C5385  ( .a(\prgm_register/n1535 ), .b(
        \prgm_register/n1536 ), .out(\prgm_register/or_signal [767]) );
  nand2 \prgm_register/C5386  ( .a(enable), .b(a[767]), .out(
        \prgm_register/n1537 ) );
  nand2 \prgm_register/C5387  ( .a(\prgm_register/en_not ), .b(a[768]), .out(
        \prgm_register/n1538 ) );
  nand2 \prgm_register/C5388  ( .a(\prgm_register/n1537 ), .b(
        \prgm_register/n1538 ), .out(\prgm_register/or_signal [768]) );
  nand2 \prgm_register/C5389  ( .a(enable), .b(a[768]), .out(
        \prgm_register/n1539 ) );
  nand2 \prgm_register/C5390  ( .a(\prgm_register/en_not ), .b(a[769]), .out(
        \prgm_register/n1540 ) );
  nand2 \prgm_register/C5391  ( .a(\prgm_register/n1539 ), .b(
        \prgm_register/n1540 ), .out(\prgm_register/or_signal [769]) );
  nand2 \prgm_register/C5392  ( .a(enable), .b(a[769]), .out(
        \prgm_register/n1541 ) );
  nand2 \prgm_register/C5393  ( .a(\prgm_register/en_not ), .b(a[770]), .out(
        \prgm_register/n1542 ) );
  nand2 \prgm_register/C5394  ( .a(\prgm_register/n1541 ), .b(
        \prgm_register/n1542 ), .out(\prgm_register/or_signal [770]) );
  nand2 \prgm_register/C5395  ( .a(enable), .b(a[770]), .out(
        \prgm_register/n1543 ) );
  nand2 \prgm_register/C5396  ( .a(\prgm_register/en_not ), .b(a[771]), .out(
        \prgm_register/n1544 ) );
  nand2 \prgm_register/C5397  ( .a(\prgm_register/n1543 ), .b(
        \prgm_register/n1544 ), .out(\prgm_register/or_signal [771]) );
  nand2 \prgm_register/C5398  ( .a(enable), .b(a[771]), .out(
        \prgm_register/n1545 ) );
  nand2 \prgm_register/C5399  ( .a(\prgm_register/en_not ), .b(a[772]), .out(
        \prgm_register/n1546 ) );
  nand2 \prgm_register/C5400  ( .a(\prgm_register/n1545 ), .b(
        \prgm_register/n1546 ), .out(\prgm_register/or_signal [772]) );
  nand2 \prgm_register/C5401  ( .a(enable), .b(a[772]), .out(
        \prgm_register/n1547 ) );
  nand2 \prgm_register/C5402  ( .a(\prgm_register/en_not ), .b(a[773]), .out(
        \prgm_register/n1548 ) );
  nand2 \prgm_register/C5403  ( .a(\prgm_register/n1547 ), .b(
        \prgm_register/n1548 ), .out(\prgm_register/or_signal [773]) );
  nand2 \prgm_register/C5404  ( .a(enable), .b(a[773]), .out(
        \prgm_register/n1549 ) );
  nand2 \prgm_register/C5405  ( .a(\prgm_register/en_not ), .b(a[774]), .out(
        \prgm_register/n1550 ) );
  nand2 \prgm_register/C5406  ( .a(\prgm_register/n1549 ), .b(
        \prgm_register/n1550 ), .out(\prgm_register/or_signal [774]) );
  nand2 \prgm_register/C5407  ( .a(enable), .b(a[774]), .out(
        \prgm_register/n1551 ) );
  nand2 \prgm_register/C5408  ( .a(\prgm_register/en_not ), .b(a[775]), .out(
        \prgm_register/n1552 ) );
  nand2 \prgm_register/C5409  ( .a(\prgm_register/n1551 ), .b(
        \prgm_register/n1552 ), .out(\prgm_register/or_signal [775]) );
  nand2 \prgm_register/C5410  ( .a(enable), .b(a[775]), .out(
        \prgm_register/n1553 ) );
  nand2 \prgm_register/C5411  ( .a(\prgm_register/en_not ), .b(a[776]), .out(
        \prgm_register/n1554 ) );
  nand2 \prgm_register/C5412  ( .a(\prgm_register/n1553 ), .b(
        \prgm_register/n1554 ), .out(\prgm_register/or_signal [776]) );
  nand2 \prgm_register/C5413  ( .a(enable), .b(a[776]), .out(
        \prgm_register/n1555 ) );
  nand2 \prgm_register/C5414  ( .a(\prgm_register/en_not ), .b(a[777]), .out(
        \prgm_register/n1556 ) );
  nand2 \prgm_register/C5415  ( .a(\prgm_register/n1555 ), .b(
        \prgm_register/n1556 ), .out(\prgm_register/or_signal [777]) );
  nand2 \prgm_register/C5416  ( .a(enable), .b(a[777]), .out(
        \prgm_register/n1557 ) );
  nand2 \prgm_register/C5417  ( .a(\prgm_register/en_not ), .b(a[778]), .out(
        \prgm_register/n1558 ) );
  nand2 \prgm_register/C5418  ( .a(\prgm_register/n1557 ), .b(
        \prgm_register/n1558 ), .out(\prgm_register/or_signal [778]) );
  nand2 \prgm_register/C5419  ( .a(enable), .b(a[778]), .out(
        \prgm_register/n1559 ) );
  nand2 \prgm_register/C5420  ( .a(\prgm_register/en_not ), .b(a[779]), .out(
        \prgm_register/n1560 ) );
  nand2 \prgm_register/C5421  ( .a(\prgm_register/n1559 ), .b(
        \prgm_register/n1560 ), .out(\prgm_register/or_signal [779]) );
  nand2 \prgm_register/C5422  ( .a(enable), .b(a[779]), .out(
        \prgm_register/n1561 ) );
  nand2 \prgm_register/C5423  ( .a(\prgm_register/en_not ), .b(a[780]), .out(
        \prgm_register/n1562 ) );
  nand2 \prgm_register/C5424  ( .a(\prgm_register/n1561 ), .b(
        \prgm_register/n1562 ), .out(\prgm_register/or_signal [780]) );
  nand2 \prgm_register/C5425  ( .a(enable), .b(a[780]), .out(
        \prgm_register/n1563 ) );
  nand2 \prgm_register/C5426  ( .a(\prgm_register/en_not ), .b(a[781]), .out(
        \prgm_register/n1564 ) );
  nand2 \prgm_register/C5427  ( .a(\prgm_register/n1563 ), .b(
        \prgm_register/n1564 ), .out(\prgm_register/or_signal [781]) );
  nand2 \prgm_register/C5428  ( .a(enable), .b(a[781]), .out(
        \prgm_register/n1565 ) );
  nand2 \prgm_register/C5429  ( .a(\prgm_register/en_not ), .b(a[782]), .out(
        \prgm_register/n1566 ) );
  nand2 \prgm_register/C5430  ( .a(\prgm_register/n1565 ), .b(
        \prgm_register/n1566 ), .out(\prgm_register/or_signal [782]) );
  nand2 \prgm_register/C5431  ( .a(enable), .b(a[782]), .out(
        \prgm_register/n1567 ) );
  nand2 \prgm_register/C5432  ( .a(\prgm_register/en_not ), .b(a[783]), .out(
        \prgm_register/n1568 ) );
  nand2 \prgm_register/C5433  ( .a(\prgm_register/n1567 ), .b(
        \prgm_register/n1568 ), .out(\prgm_register/or_signal [783]) );
  nand2 \prgm_register/C5434  ( .a(enable), .b(a[783]), .out(
        \prgm_register/n1569 ) );
  nand2 \prgm_register/C5435  ( .a(\prgm_register/en_not ), .b(a[784]), .out(
        \prgm_register/n1570 ) );
  nand2 \prgm_register/C5436  ( .a(\prgm_register/n1569 ), .b(
        \prgm_register/n1570 ), .out(\prgm_register/or_signal [784]) );
  nand2 \prgm_register/C5437  ( .a(enable), .b(a[784]), .out(
        \prgm_register/n1571 ) );
  nand2 \prgm_register/C5438  ( .a(\prgm_register/en_not ), .b(a[785]), .out(
        \prgm_register/n1572 ) );
  nand2 \prgm_register/C5439  ( .a(\prgm_register/n1571 ), .b(
        \prgm_register/n1572 ), .out(\prgm_register/or_signal [785]) );
  nand2 \prgm_register/C5440  ( .a(enable), .b(a[785]), .out(
        \prgm_register/n1573 ) );
  nand2 \prgm_register/C5441  ( .a(\prgm_register/en_not ), .b(a[786]), .out(
        \prgm_register/n1574 ) );
  nand2 \prgm_register/C5442  ( .a(\prgm_register/n1573 ), .b(
        \prgm_register/n1574 ), .out(\prgm_register/or_signal [786]) );
  nand2 \prgm_register/C5443  ( .a(enable), .b(a[786]), .out(
        \prgm_register/n1575 ) );
  nand2 \prgm_register/C5444  ( .a(\prgm_register/en_not ), .b(a[787]), .out(
        \prgm_register/n1576 ) );
  nand2 \prgm_register/C5445  ( .a(\prgm_register/n1575 ), .b(
        \prgm_register/n1576 ), .out(\prgm_register/or_signal [787]) );
  nand2 \prgm_register/C5446  ( .a(enable), .b(a[787]), .out(
        \prgm_register/n1577 ) );
  nand2 \prgm_register/C5447  ( .a(\prgm_register/en_not ), .b(a[788]), .out(
        \prgm_register/n1578 ) );
  nand2 \prgm_register/C5448  ( .a(\prgm_register/n1577 ), .b(
        \prgm_register/n1578 ), .out(\prgm_register/or_signal [788]) );
  nand2 \prgm_register/C5449  ( .a(enable), .b(a[788]), .out(
        \prgm_register/n1579 ) );
  nand2 \prgm_register/C5450  ( .a(\prgm_register/en_not ), .b(a[789]), .out(
        \prgm_register/n1580 ) );
  nand2 \prgm_register/C5451  ( .a(\prgm_register/n1579 ), .b(
        \prgm_register/n1580 ), .out(\prgm_register/or_signal [789]) );
  nand2 \prgm_register/C5452  ( .a(enable), .b(a[789]), .out(
        \prgm_register/n1581 ) );
  nand2 \prgm_register/C5453  ( .a(\prgm_register/en_not ), .b(a[790]), .out(
        \prgm_register/n1582 ) );
  nand2 \prgm_register/C5454  ( .a(\prgm_register/n1581 ), .b(
        \prgm_register/n1582 ), .out(\prgm_register/or_signal [790]) );
  nand2 \prgm_register/C5455  ( .a(enable), .b(a[790]), .out(
        \prgm_register/n1583 ) );
  nand2 \prgm_register/C5456  ( .a(\prgm_register/en_not ), .b(a[791]), .out(
        \prgm_register/n1584 ) );
  nand2 \prgm_register/C5457  ( .a(\prgm_register/n1583 ), .b(
        \prgm_register/n1584 ), .out(\prgm_register/or_signal [791]) );
  nand2 \prgm_register/C5458  ( .a(enable), .b(a[791]), .out(
        \prgm_register/n1585 ) );
  nand2 \prgm_register/C5459  ( .a(\prgm_register/en_not ), .b(a[792]), .out(
        \prgm_register/n1586 ) );
  nand2 \prgm_register/C5460  ( .a(\prgm_register/n1585 ), .b(
        \prgm_register/n1586 ), .out(\prgm_register/or_signal [792]) );
  nand2 \prgm_register/C5461  ( .a(enable), .b(a[792]), .out(
        \prgm_register/n1587 ) );
  nand2 \prgm_register/C5462  ( .a(\prgm_register/en_not ), .b(a[793]), .out(
        \prgm_register/n1588 ) );
  nand2 \prgm_register/C5463  ( .a(\prgm_register/n1587 ), .b(
        \prgm_register/n1588 ), .out(\prgm_register/or_signal [793]) );
  nand2 \prgm_register/C5464  ( .a(enable), .b(a[793]), .out(
        \prgm_register/n1589 ) );
  nand2 \prgm_register/C5465  ( .a(\prgm_register/en_not ), .b(a[794]), .out(
        \prgm_register/n1590 ) );
  nand2 \prgm_register/C5466  ( .a(\prgm_register/n1589 ), .b(
        \prgm_register/n1590 ), .out(\prgm_register/or_signal [794]) );
  nand2 \prgm_register/C5467  ( .a(enable), .b(a[794]), .out(
        \prgm_register/n1591 ) );
  nand2 \prgm_register/C5468  ( .a(\prgm_register/en_not ), .b(a[795]), .out(
        \prgm_register/n1592 ) );
  nand2 \prgm_register/C5469  ( .a(\prgm_register/n1591 ), .b(
        \prgm_register/n1592 ), .out(\prgm_register/or_signal [795]) );
  nand2 \prgm_register/C5470  ( .a(enable), .b(a[795]), .out(
        \prgm_register/n1593 ) );
  nand2 \prgm_register/C5471  ( .a(\prgm_register/en_not ), .b(a[796]), .out(
        \prgm_register/n1594 ) );
  nand2 \prgm_register/C5472  ( .a(\prgm_register/n1593 ), .b(
        \prgm_register/n1594 ), .out(\prgm_register/or_signal [796]) );
  nand2 \prgm_register/C5473  ( .a(enable), .b(a[796]), .out(
        \prgm_register/n1595 ) );
  nand2 \prgm_register/C5474  ( .a(\prgm_register/en_not ), .b(a[797]), .out(
        \prgm_register/n1596 ) );
  nand2 \prgm_register/C5475  ( .a(\prgm_register/n1595 ), .b(
        \prgm_register/n1596 ), .out(\prgm_register/or_signal [797]) );
  nand2 \prgm_register/C5476  ( .a(enable), .b(a[797]), .out(
        \prgm_register/n1597 ) );
  nand2 \prgm_register/C5477  ( .a(\prgm_register/en_not ), .b(a[798]), .out(
        \prgm_register/n1598 ) );
  nand2 \prgm_register/C5478  ( .a(\prgm_register/n1597 ), .b(
        \prgm_register/n1598 ), .out(\prgm_register/or_signal [798]) );
  nand2 \prgm_register/C5479  ( .a(enable), .b(a[798]), .out(
        \prgm_register/n1599 ) );
  nand2 \prgm_register/C5480  ( .a(\prgm_register/en_not ), .b(a[799]), .out(
        \prgm_register/n1600 ) );
  nand2 \prgm_register/C5481  ( .a(\prgm_register/n1599 ), .b(
        \prgm_register/n1600 ), .out(\prgm_register/or_signal [799]) );
  nand2 \prgm_register/C5482  ( .a(enable), .b(a[799]), .out(
        \prgm_register/n1601 ) );
  nand2 \prgm_register/C5483  ( .a(\prgm_register/en_not ), .b(a[800]), .out(
        \prgm_register/n1602 ) );
  nand2 \prgm_register/C5484  ( .a(\prgm_register/n1601 ), .b(
        \prgm_register/n1602 ), .out(\prgm_register/or_signal [800]) );
  nand2 \prgm_register/C5485  ( .a(enable), .b(a[800]), .out(
        \prgm_register/n1603 ) );
  nand2 \prgm_register/C5486  ( .a(\prgm_register/en_not ), .b(a[801]), .out(
        \prgm_register/n1604 ) );
  nand2 \prgm_register/C5487  ( .a(\prgm_register/n1603 ), .b(
        \prgm_register/n1604 ), .out(\prgm_register/or_signal [801]) );
  nand2 \prgm_register/C5488  ( .a(enable), .b(a[801]), .out(
        \prgm_register/n1605 ) );
  nand2 \prgm_register/C5489  ( .a(\prgm_register/en_not ), .b(a[802]), .out(
        \prgm_register/n1606 ) );
  nand2 \prgm_register/C5490  ( .a(\prgm_register/n1605 ), .b(
        \prgm_register/n1606 ), .out(\prgm_register/or_signal [802]) );
  nand2 \prgm_register/C5491  ( .a(enable), .b(a[802]), .out(
        \prgm_register/n1607 ) );
  nand2 \prgm_register/C5492  ( .a(\prgm_register/en_not ), .b(a[803]), .out(
        \prgm_register/n1608 ) );
  nand2 \prgm_register/C5493  ( .a(\prgm_register/n1607 ), .b(
        \prgm_register/n1608 ), .out(\prgm_register/or_signal [803]) );
  nand2 \prgm_register/C5494  ( .a(enable), .b(a[803]), .out(
        \prgm_register/n1609 ) );
  nand2 \prgm_register/C5495  ( .a(\prgm_register/en_not ), .b(a[804]), .out(
        \prgm_register/n1610 ) );
  nand2 \prgm_register/C5496  ( .a(\prgm_register/n1609 ), .b(
        \prgm_register/n1610 ), .out(\prgm_register/or_signal [804]) );
  nand2 \prgm_register/C5497  ( .a(enable), .b(a[804]), .out(
        \prgm_register/n1611 ) );
  nand2 \prgm_register/C5498  ( .a(\prgm_register/en_not ), .b(a[805]), .out(
        \prgm_register/n1612 ) );
  nand2 \prgm_register/C5499  ( .a(\prgm_register/n1611 ), .b(
        \prgm_register/n1612 ), .out(\prgm_register/or_signal [805]) );
  nand2 \prgm_register/C5500  ( .a(enable), .b(a[805]), .out(
        \prgm_register/n1613 ) );
  nand2 \prgm_register/C5501  ( .a(\prgm_register/en_not ), .b(a[806]), .out(
        \prgm_register/n1614 ) );
  nand2 \prgm_register/C5502  ( .a(\prgm_register/n1613 ), .b(
        \prgm_register/n1614 ), .out(\prgm_register/or_signal [806]) );
  nand2 \prgm_register/C5503  ( .a(enable), .b(a[806]), .out(
        \prgm_register/n1615 ) );
  nand2 \prgm_register/C5504  ( .a(\prgm_register/en_not ), .b(a[807]), .out(
        \prgm_register/n1616 ) );
  nand2 \prgm_register/C5505  ( .a(\prgm_register/n1615 ), .b(
        \prgm_register/n1616 ), .out(\prgm_register/or_signal [807]) );
  nand2 \prgm_register/C5506  ( .a(enable), .b(a[807]), .out(
        \prgm_register/n1617 ) );
  nand2 \prgm_register/C5507  ( .a(\prgm_register/en_not ), .b(a[808]), .out(
        \prgm_register/n1618 ) );
  nand2 \prgm_register/C5508  ( .a(\prgm_register/n1617 ), .b(
        \prgm_register/n1618 ), .out(\prgm_register/or_signal [808]) );
  nand2 \prgm_register/C5509  ( .a(enable), .b(a[808]), .out(
        \prgm_register/n1619 ) );
  nand2 \prgm_register/C5510  ( .a(\prgm_register/en_not ), .b(a[809]), .out(
        \prgm_register/n1620 ) );
  nand2 \prgm_register/C5511  ( .a(\prgm_register/n1619 ), .b(
        \prgm_register/n1620 ), .out(\prgm_register/or_signal [809]) );
  nand2 \prgm_register/C5512  ( .a(enable), .b(a[809]), .out(
        \prgm_register/n1621 ) );
  nand2 \prgm_register/C5513  ( .a(\prgm_register/en_not ), .b(a[810]), .out(
        \prgm_register/n1622 ) );
  nand2 \prgm_register/C5514  ( .a(\prgm_register/n1621 ), .b(
        \prgm_register/n1622 ), .out(\prgm_register/or_signal [810]) );
  nand2 \prgm_register/C5515  ( .a(enable), .b(a[810]), .out(
        \prgm_register/n1623 ) );
  nand2 \prgm_register/C5516  ( .a(\prgm_register/en_not ), .b(a[811]), .out(
        \prgm_register/n1624 ) );
  nand2 \prgm_register/C5517  ( .a(\prgm_register/n1623 ), .b(
        \prgm_register/n1624 ), .out(\prgm_register/or_signal [811]) );
  nand2 \prgm_register/C5518  ( .a(enable), .b(a[811]), .out(
        \prgm_register/n1625 ) );
  nand2 \prgm_register/C5519  ( .a(\prgm_register/en_not ), .b(a[812]), .out(
        \prgm_register/n1626 ) );
  nand2 \prgm_register/C5520  ( .a(\prgm_register/n1625 ), .b(
        \prgm_register/n1626 ), .out(\prgm_register/or_signal [812]) );
  nand2 \prgm_register/C5521  ( .a(enable), .b(a[812]), .out(
        \prgm_register/n1627 ) );
  nand2 \prgm_register/C5522  ( .a(\prgm_register/en_not ), .b(a[813]), .out(
        \prgm_register/n1628 ) );
  nand2 \prgm_register/C5523  ( .a(\prgm_register/n1627 ), .b(
        \prgm_register/n1628 ), .out(\prgm_register/or_signal [813]) );
  nand2 \prgm_register/C5524  ( .a(enable), .b(a[813]), .out(
        \prgm_register/n1629 ) );
  nand2 \prgm_register/C5525  ( .a(\prgm_register/en_not ), .b(a[814]), .out(
        \prgm_register/n1630 ) );
  nand2 \prgm_register/C5526  ( .a(\prgm_register/n1629 ), .b(
        \prgm_register/n1630 ), .out(\prgm_register/or_signal [814]) );
  nand2 \prgm_register/C5527  ( .a(enable), .b(a[814]), .out(
        \prgm_register/n1631 ) );
  nand2 \prgm_register/C5528  ( .a(\prgm_register/en_not ), .b(a[815]), .out(
        \prgm_register/n1632 ) );
  nand2 \prgm_register/C5529  ( .a(\prgm_register/n1631 ), .b(
        \prgm_register/n1632 ), .out(\prgm_register/or_signal [815]) );
  nand2 \prgm_register/C5530  ( .a(enable), .b(a[815]), .out(
        \prgm_register/n1633 ) );
  nand2 \prgm_register/C5531  ( .a(\prgm_register/en_not ), .b(a[816]), .out(
        \prgm_register/n1634 ) );
  nand2 \prgm_register/C5532  ( .a(\prgm_register/n1633 ), .b(
        \prgm_register/n1634 ), .out(\prgm_register/or_signal [816]) );
  nand2 \prgm_register/C5533  ( .a(enable), .b(a[816]), .out(
        \prgm_register/n1635 ) );
  nand2 \prgm_register/C5534  ( .a(\prgm_register/en_not ), .b(a[817]), .out(
        \prgm_register/n1636 ) );
  nand2 \prgm_register/C5535  ( .a(\prgm_register/n1635 ), .b(
        \prgm_register/n1636 ), .out(\prgm_register/or_signal [817]) );
  nand2 \prgm_register/C5536  ( .a(enable), .b(a[817]), .out(
        \prgm_register/n1637 ) );
  nand2 \prgm_register/C5537  ( .a(\prgm_register/en_not ), .b(a[818]), .out(
        \prgm_register/n1638 ) );
  nand2 \prgm_register/C5538  ( .a(\prgm_register/n1637 ), .b(
        \prgm_register/n1638 ), .out(\prgm_register/or_signal [818]) );
  nand2 \prgm_register/C5539  ( .a(enable), .b(a[818]), .out(
        \prgm_register/n1639 ) );
  nand2 \prgm_register/C5540  ( .a(\prgm_register/en_not ), .b(a[819]), .out(
        \prgm_register/n1640 ) );
  nand2 \prgm_register/C5541  ( .a(\prgm_register/n1639 ), .b(
        \prgm_register/n1640 ), .out(\prgm_register/or_signal [819]) );
  nand2 \prgm_register/C5542  ( .a(enable), .b(a[819]), .out(
        \prgm_register/n1641 ) );
  nand2 \prgm_register/C5543  ( .a(\prgm_register/en_not ), .b(a[820]), .out(
        \prgm_register/n1642 ) );
  nand2 \prgm_register/C5544  ( .a(\prgm_register/n1641 ), .b(
        \prgm_register/n1642 ), .out(\prgm_register/or_signal [820]) );
  nand2 \prgm_register/C5545  ( .a(enable), .b(a[820]), .out(
        \prgm_register/n1643 ) );
  nand2 \prgm_register/C5546  ( .a(\prgm_register/en_not ), .b(a[821]), .out(
        \prgm_register/n1644 ) );
  nand2 \prgm_register/C5547  ( .a(\prgm_register/n1643 ), .b(
        \prgm_register/n1644 ), .out(\prgm_register/or_signal [821]) );
  nand2 \prgm_register/C5548  ( .a(enable), .b(a[821]), .out(
        \prgm_register/n1645 ) );
  nand2 \prgm_register/C5549  ( .a(\prgm_register/en_not ), .b(a[822]), .out(
        \prgm_register/n1646 ) );
  nand2 \prgm_register/C5550  ( .a(\prgm_register/n1645 ), .b(
        \prgm_register/n1646 ), .out(\prgm_register/or_signal [822]) );
  nand2 \prgm_register/C5551  ( .a(enable), .b(a[822]), .out(
        \prgm_register/n1647 ) );
  nand2 \prgm_register/C5552  ( .a(\prgm_register/en_not ), .b(a[823]), .out(
        \prgm_register/n1648 ) );
  nand2 \prgm_register/C5553  ( .a(\prgm_register/n1647 ), .b(
        \prgm_register/n1648 ), .out(\prgm_register/or_signal [823]) );
  nand2 \prgm_register/C5554  ( .a(enable), .b(a[823]), .out(
        \prgm_register/n1649 ) );
  nand2 \prgm_register/C5555  ( .a(\prgm_register/en_not ), .b(a[824]), .out(
        \prgm_register/n1650 ) );
  nand2 \prgm_register/C5556  ( .a(\prgm_register/n1649 ), .b(
        \prgm_register/n1650 ), .out(\prgm_register/or_signal [824]) );
  nand2 \prgm_register/C5557  ( .a(enable), .b(a[824]), .out(
        \prgm_register/n1651 ) );
  nand2 \prgm_register/C5558  ( .a(\prgm_register/en_not ), .b(a[825]), .out(
        \prgm_register/n1652 ) );
  nand2 \prgm_register/C5559  ( .a(\prgm_register/n1651 ), .b(
        \prgm_register/n1652 ), .out(\prgm_register/or_signal [825]) );
  nand2 \prgm_register/C5560  ( .a(enable), .b(a[825]), .out(
        \prgm_register/n1653 ) );
  nand2 \prgm_register/C5561  ( .a(\prgm_register/en_not ), .b(a[826]), .out(
        \prgm_register/n1654 ) );
  nand2 \prgm_register/C5562  ( .a(\prgm_register/n1653 ), .b(
        \prgm_register/n1654 ), .out(\prgm_register/or_signal [826]) );
  nand2 \prgm_register/C5563  ( .a(enable), .b(a[826]), .out(
        \prgm_register/n1655 ) );
  nand2 \prgm_register/C5564  ( .a(\prgm_register/en_not ), .b(a[827]), .out(
        \prgm_register/n1656 ) );
  nand2 \prgm_register/C5565  ( .a(\prgm_register/n1655 ), .b(
        \prgm_register/n1656 ), .out(\prgm_register/or_signal [827]) );
  nand2 \prgm_register/C5566  ( .a(enable), .b(a[827]), .out(
        \prgm_register/n1657 ) );
  nand2 \prgm_register/C5567  ( .a(\prgm_register/en_not ), .b(a[828]), .out(
        \prgm_register/n1658 ) );
  nand2 \prgm_register/C5568  ( .a(\prgm_register/n1657 ), .b(
        \prgm_register/n1658 ), .out(\prgm_register/or_signal [828]) );
  nand2 \prgm_register/C5569  ( .a(enable), .b(a[828]), .out(
        \prgm_register/n1659 ) );
  nand2 \prgm_register/C5570  ( .a(\prgm_register/en_not ), .b(a[829]), .out(
        \prgm_register/n1660 ) );
  nand2 \prgm_register/C5571  ( .a(\prgm_register/n1659 ), .b(
        \prgm_register/n1660 ), .out(\prgm_register/or_signal [829]) );
  nand2 \prgm_register/C5572  ( .a(enable), .b(a[829]), .out(
        \prgm_register/n1661 ) );
  nand2 \prgm_register/C5573  ( .a(\prgm_register/en_not ), .b(a[830]), .out(
        \prgm_register/n1662 ) );
  nand2 \prgm_register/C5574  ( .a(\prgm_register/n1661 ), .b(
        \prgm_register/n1662 ), .out(\prgm_register/or_signal [830]) );
  nand2 \prgm_register/C5575  ( .a(enable), .b(a[830]), .out(
        \prgm_register/n1663 ) );
  nand2 \prgm_register/C5576  ( .a(\prgm_register/en_not ), .b(a[831]), .out(
        \prgm_register/n1664 ) );
  nand2 \prgm_register/C5577  ( .a(\prgm_register/n1663 ), .b(
        \prgm_register/n1664 ), .out(\prgm_register/or_signal [831]) );
  nand2 \prgm_register/C5578  ( .a(enable), .b(a[831]), .out(
        \prgm_register/n1665 ) );
  nand2 \prgm_register/C5579  ( .a(\prgm_register/en_not ), .b(a[832]), .out(
        \prgm_register/n1666 ) );
  nand2 \prgm_register/C5580  ( .a(\prgm_register/n1665 ), .b(
        \prgm_register/n1666 ), .out(\prgm_register/or_signal [832]) );
  nand2 \prgm_register/C5581  ( .a(enable), .b(a[832]), .out(
        \prgm_register/n1667 ) );
  nand2 \prgm_register/C5582  ( .a(\prgm_register/en_not ), .b(a[833]), .out(
        \prgm_register/n1668 ) );
  nand2 \prgm_register/C5583  ( .a(\prgm_register/n1667 ), .b(
        \prgm_register/n1668 ), .out(\prgm_register/or_signal [833]) );
  nand2 \prgm_register/C5584  ( .a(enable), .b(a[833]), .out(
        \prgm_register/n1669 ) );
  nand2 \prgm_register/C5585  ( .a(\prgm_register/en_not ), .b(a[834]), .out(
        \prgm_register/n1670 ) );
  nand2 \prgm_register/C5586  ( .a(\prgm_register/n1669 ), .b(
        \prgm_register/n1670 ), .out(\prgm_register/or_signal [834]) );
  nand2 \prgm_register/C5587  ( .a(enable), .b(a[834]), .out(
        \prgm_register/n1671 ) );
  nand2 \prgm_register/C5588  ( .a(\prgm_register/en_not ), .b(a[835]), .out(
        \prgm_register/n1672 ) );
  nand2 \prgm_register/C5589  ( .a(\prgm_register/n1671 ), .b(
        \prgm_register/n1672 ), .out(\prgm_register/or_signal [835]) );
  nand2 \prgm_register/C5590  ( .a(enable), .b(a[835]), .out(
        \prgm_register/n1673 ) );
  nand2 \prgm_register/C5591  ( .a(\prgm_register/en_not ), .b(a[836]), .out(
        \prgm_register/n1674 ) );
  nand2 \prgm_register/C5592  ( .a(\prgm_register/n1673 ), .b(
        \prgm_register/n1674 ), .out(\prgm_register/or_signal [836]) );
  nand2 \prgm_register/C5593  ( .a(enable), .b(a[836]), .out(
        \prgm_register/n1675 ) );
  nand2 \prgm_register/C5594  ( .a(\prgm_register/en_not ), .b(a[837]), .out(
        \prgm_register/n1676 ) );
  nand2 \prgm_register/C5595  ( .a(\prgm_register/n1675 ), .b(
        \prgm_register/n1676 ), .out(\prgm_register/or_signal [837]) );
  nand2 \prgm_register/C5596  ( .a(enable), .b(a[837]), .out(
        \prgm_register/n1677 ) );
  nand2 \prgm_register/C5597  ( .a(\prgm_register/en_not ), .b(a[838]), .out(
        \prgm_register/n1678 ) );
  nand2 \prgm_register/C5598  ( .a(\prgm_register/n1677 ), .b(
        \prgm_register/n1678 ), .out(\prgm_register/or_signal [838]) );
  nand2 \prgm_register/C5599  ( .a(enable), .b(a[838]), .out(
        \prgm_register/n1679 ) );
  nand2 \prgm_register/C5600  ( .a(\prgm_register/en_not ), .b(a[839]), .out(
        \prgm_register/n1680 ) );
  nand2 \prgm_register/C5601  ( .a(\prgm_register/n1679 ), .b(
        \prgm_register/n1680 ), .out(\prgm_register/or_signal [839]) );
  nand2 \prgm_register/C5602  ( .a(enable), .b(a[839]), .out(
        \prgm_register/n1681 ) );
  nand2 \prgm_register/C5603  ( .a(\prgm_register/en_not ), .b(a[840]), .out(
        \prgm_register/n1682 ) );
  nand2 \prgm_register/C5604  ( .a(\prgm_register/n1681 ), .b(
        \prgm_register/n1682 ), .out(\prgm_register/or_signal [840]) );
  nand2 \prgm_register/C5605  ( .a(enable), .b(a[840]), .out(
        \prgm_register/n1683 ) );
  nand2 \prgm_register/C5606  ( .a(\prgm_register/en_not ), .b(a[841]), .out(
        \prgm_register/n1684 ) );
  nand2 \prgm_register/C5607  ( .a(\prgm_register/n1683 ), .b(
        \prgm_register/n1684 ), .out(\prgm_register/or_signal [841]) );
  nand2 \prgm_register/C5608  ( .a(enable), .b(a[841]), .out(
        \prgm_register/n1685 ) );
  nand2 \prgm_register/C5609  ( .a(\prgm_register/en_not ), .b(a[842]), .out(
        \prgm_register/n1686 ) );
  nand2 \prgm_register/C5610  ( .a(\prgm_register/n1685 ), .b(
        \prgm_register/n1686 ), .out(\prgm_register/or_signal [842]) );
  nand2 \prgm_register/C5611  ( .a(enable), .b(a[842]), .out(
        \prgm_register/n1687 ) );
  nand2 \prgm_register/C5612  ( .a(\prgm_register/en_not ), .b(a[843]), .out(
        \prgm_register/n1688 ) );
  nand2 \prgm_register/C5613  ( .a(\prgm_register/n1687 ), .b(
        \prgm_register/n1688 ), .out(\prgm_register/or_signal [843]) );
  nand2 \prgm_register/C5614  ( .a(enable), .b(a[843]), .out(
        \prgm_register/n1689 ) );
  nand2 \prgm_register/C5615  ( .a(\prgm_register/en_not ), .b(a[844]), .out(
        \prgm_register/n1690 ) );
  nand2 \prgm_register/C5616  ( .a(\prgm_register/n1689 ), .b(
        \prgm_register/n1690 ), .out(\prgm_register/or_signal [844]) );
  nand2 \prgm_register/C5617  ( .a(enable), .b(a[844]), .out(
        \prgm_register/n1691 ) );
  nand2 \prgm_register/C5618  ( .a(\prgm_register/en_not ), .b(a[845]), .out(
        \prgm_register/n1692 ) );
  nand2 \prgm_register/C5619  ( .a(\prgm_register/n1691 ), .b(
        \prgm_register/n1692 ), .out(\prgm_register/or_signal [845]) );
  nand2 \prgm_register/C5620  ( .a(enable), .b(a[845]), .out(
        \prgm_register/n1693 ) );
  nand2 \prgm_register/C5621  ( .a(\prgm_register/en_not ), .b(a[846]), .out(
        \prgm_register/n1694 ) );
  nand2 \prgm_register/C5622  ( .a(\prgm_register/n1693 ), .b(
        \prgm_register/n1694 ), .out(\prgm_register/or_signal [846]) );
  nand2 \prgm_register/C5623  ( .a(enable), .b(a[846]), .out(
        \prgm_register/n1695 ) );
  nand2 \prgm_register/C5624  ( .a(\prgm_register/en_not ), .b(a[847]), .out(
        \prgm_register/n1696 ) );
  nand2 \prgm_register/C5625  ( .a(\prgm_register/n1695 ), .b(
        \prgm_register/n1696 ), .out(\prgm_register/or_signal [847]) );
  nand2 \prgm_register/C5626  ( .a(enable), .b(a[847]), .out(
        \prgm_register/n1697 ) );
  nand2 \prgm_register/C5627  ( .a(\prgm_register/en_not ), .b(a[848]), .out(
        \prgm_register/n1698 ) );
  nand2 \prgm_register/C5628  ( .a(\prgm_register/n1697 ), .b(
        \prgm_register/n1698 ), .out(\prgm_register/or_signal [848]) );
  nand2 \prgm_register/C5629  ( .a(enable), .b(a[848]), .out(
        \prgm_register/n1699 ) );
  nand2 \prgm_register/C5630  ( .a(\prgm_register/en_not ), .b(a[849]), .out(
        \prgm_register/n1700 ) );
  nand2 \prgm_register/C5631  ( .a(\prgm_register/n1699 ), .b(
        \prgm_register/n1700 ), .out(\prgm_register/or_signal [849]) );
  nand2 \prgm_register/C5632  ( .a(enable), .b(a[849]), .out(
        \prgm_register/n1701 ) );
  nand2 \prgm_register/C5633  ( .a(\prgm_register/en_not ), .b(a[850]), .out(
        \prgm_register/n1702 ) );
  nand2 \prgm_register/C5634  ( .a(\prgm_register/n1701 ), .b(
        \prgm_register/n1702 ), .out(\prgm_register/or_signal [850]) );
  nand2 \prgm_register/C5635  ( .a(enable), .b(a[850]), .out(
        \prgm_register/n1703 ) );
  nand2 \prgm_register/C5636  ( .a(\prgm_register/en_not ), .b(a[851]), .out(
        \prgm_register/n1704 ) );
  nand2 \prgm_register/C5637  ( .a(\prgm_register/n1703 ), .b(
        \prgm_register/n1704 ), .out(\prgm_register/or_signal [851]) );
  nand2 \prgm_register/C5638  ( .a(enable), .b(a[851]), .out(
        \prgm_register/n1705 ) );
  nand2 \prgm_register/C5639  ( .a(\prgm_register/en_not ), .b(a[852]), .out(
        \prgm_register/n1706 ) );
  nand2 \prgm_register/C5640  ( .a(\prgm_register/n1705 ), .b(
        \prgm_register/n1706 ), .out(\prgm_register/or_signal [852]) );
  nand2 \prgm_register/C5641  ( .a(enable), .b(a[852]), .out(
        \prgm_register/n1707 ) );
  nand2 \prgm_register/C5642  ( .a(\prgm_register/en_not ), .b(a[853]), .out(
        \prgm_register/n1708 ) );
  nand2 \prgm_register/C5643  ( .a(\prgm_register/n1707 ), .b(
        \prgm_register/n1708 ), .out(\prgm_register/or_signal [853]) );
  nand2 \prgm_register/C5644  ( .a(enable), .b(a[853]), .out(
        \prgm_register/n1709 ) );
  nand2 \prgm_register/C5645  ( .a(\prgm_register/en_not ), .b(a[854]), .out(
        \prgm_register/n1710 ) );
  nand2 \prgm_register/C5646  ( .a(\prgm_register/n1709 ), .b(
        \prgm_register/n1710 ), .out(\prgm_register/or_signal [854]) );
  nand2 \prgm_register/C5647  ( .a(enable), .b(a[854]), .out(
        \prgm_register/n1711 ) );
  nand2 \prgm_register/C5648  ( .a(\prgm_register/en_not ), .b(a[855]), .out(
        \prgm_register/n1712 ) );
  nand2 \prgm_register/C5649  ( .a(\prgm_register/n1711 ), .b(
        \prgm_register/n1712 ), .out(\prgm_register/or_signal [855]) );
  nand2 \prgm_register/C5650  ( .a(enable), .b(a[855]), .out(
        \prgm_register/n1713 ) );
  nand2 \prgm_register/C5651  ( .a(\prgm_register/en_not ), .b(a[856]), .out(
        \prgm_register/n1714 ) );
  nand2 \prgm_register/C5652  ( .a(\prgm_register/n1713 ), .b(
        \prgm_register/n1714 ), .out(\prgm_register/or_signal [856]) );
  nand2 \prgm_register/C5653  ( .a(enable), .b(a[856]), .out(
        \prgm_register/n1715 ) );
  nand2 \prgm_register/C5654  ( .a(\prgm_register/en_not ), .b(a[857]), .out(
        \prgm_register/n1716 ) );
  nand2 \prgm_register/C5655  ( .a(\prgm_register/n1715 ), .b(
        \prgm_register/n1716 ), .out(\prgm_register/or_signal [857]) );
  nand2 \prgm_register/C5656  ( .a(enable), .b(a[857]), .out(
        \prgm_register/n1717 ) );
  nand2 \prgm_register/C5657  ( .a(\prgm_register/en_not ), .b(a[858]), .out(
        \prgm_register/n1718 ) );
  nand2 \prgm_register/C5658  ( .a(\prgm_register/n1717 ), .b(
        \prgm_register/n1718 ), .out(\prgm_register/or_signal [858]) );
  nand2 \prgm_register/C5659  ( .a(enable), .b(a[858]), .out(
        \prgm_register/n1719 ) );
  nand2 \prgm_register/C5660  ( .a(\prgm_register/en_not ), .b(a[859]), .out(
        \prgm_register/n1720 ) );
  nand2 \prgm_register/C5661  ( .a(\prgm_register/n1719 ), .b(
        \prgm_register/n1720 ), .out(\prgm_register/or_signal [859]) );
  nand2 \prgm_register/C5662  ( .a(enable), .b(a[859]), .out(
        \prgm_register/n1721 ) );
  nand2 \prgm_register/C5663  ( .a(\prgm_register/en_not ), .b(a[860]), .out(
        \prgm_register/n1722 ) );
  nand2 \prgm_register/C5664  ( .a(\prgm_register/n1721 ), .b(
        \prgm_register/n1722 ), .out(\prgm_register/or_signal [860]) );
  nand2 \prgm_register/C5665  ( .a(enable), .b(a[860]), .out(
        \prgm_register/n1723 ) );
  nand2 \prgm_register/C5666  ( .a(\prgm_register/en_not ), .b(a[861]), .out(
        \prgm_register/n1724 ) );
  nand2 \prgm_register/C5667  ( .a(\prgm_register/n1723 ), .b(
        \prgm_register/n1724 ), .out(\prgm_register/or_signal [861]) );
  nand2 \prgm_register/C5668  ( .a(enable), .b(a[861]), .out(
        \prgm_register/n1725 ) );
  nand2 \prgm_register/C5669  ( .a(\prgm_register/en_not ), .b(a[862]), .out(
        \prgm_register/n1726 ) );
  nand2 \prgm_register/C5670  ( .a(\prgm_register/n1725 ), .b(
        \prgm_register/n1726 ), .out(\prgm_register/or_signal [862]) );
  nand2 \prgm_register/C5671  ( .a(enable), .b(a[862]), .out(
        \prgm_register/n1727 ) );
  nand2 \prgm_register/C5672  ( .a(\prgm_register/en_not ), .b(a[863]), .out(
        \prgm_register/n1728 ) );
  nand2 \prgm_register/C5673  ( .a(\prgm_register/n1727 ), .b(
        \prgm_register/n1728 ), .out(\prgm_register/or_signal [863]) );
  nand2 \prgm_register/C5674  ( .a(enable), .b(a[863]), .out(
        \prgm_register/n1729 ) );
  nand2 \prgm_register/C5675  ( .a(\prgm_register/en_not ), .b(a[864]), .out(
        \prgm_register/n1730 ) );
  nand2 \prgm_register/C5676  ( .a(\prgm_register/n1729 ), .b(
        \prgm_register/n1730 ), .out(\prgm_register/or_signal [864]) );
  nand2 \prgm_register/C5677  ( .a(enable), .b(a[864]), .out(
        \prgm_register/n1731 ) );
  nand2 \prgm_register/C5678  ( .a(\prgm_register/en_not ), .b(a[865]), .out(
        \prgm_register/n1732 ) );
  nand2 \prgm_register/C5679  ( .a(\prgm_register/n1731 ), .b(
        \prgm_register/n1732 ), .out(\prgm_register/or_signal [865]) );
  nand2 \prgm_register/C5680  ( .a(enable), .b(a[865]), .out(
        \prgm_register/n1733 ) );
  nand2 \prgm_register/C5681  ( .a(\prgm_register/en_not ), .b(a[866]), .out(
        \prgm_register/n1734 ) );
  nand2 \prgm_register/C5682  ( .a(\prgm_register/n1733 ), .b(
        \prgm_register/n1734 ), .out(\prgm_register/or_signal [866]) );
  nand2 \prgm_register/C5683  ( .a(enable), .b(a[866]), .out(
        \prgm_register/n1735 ) );
  nand2 \prgm_register/C5684  ( .a(\prgm_register/en_not ), .b(a[867]), .out(
        \prgm_register/n1736 ) );
  nand2 \prgm_register/C5685  ( .a(\prgm_register/n1735 ), .b(
        \prgm_register/n1736 ), .out(\prgm_register/or_signal [867]) );
  nand2 \prgm_register/C5686  ( .a(enable), .b(a[867]), .out(
        \prgm_register/n1737 ) );
  nand2 \prgm_register/C5687  ( .a(\prgm_register/en_not ), .b(a[868]), .out(
        \prgm_register/n1738 ) );
  nand2 \prgm_register/C5688  ( .a(\prgm_register/n1737 ), .b(
        \prgm_register/n1738 ), .out(\prgm_register/or_signal [868]) );
  nand2 \prgm_register/C5689  ( .a(enable), .b(a[868]), .out(
        \prgm_register/n1739 ) );
  nand2 \prgm_register/C5690  ( .a(\prgm_register/en_not ), .b(a[869]), .out(
        \prgm_register/n1740 ) );
  nand2 \prgm_register/C5691  ( .a(\prgm_register/n1739 ), .b(
        \prgm_register/n1740 ), .out(\prgm_register/or_signal [869]) );
  nand2 \prgm_register/C5692  ( .a(enable), .b(a[869]), .out(
        \prgm_register/n1741 ) );
  nand2 \prgm_register/C5693  ( .a(\prgm_register/en_not ), .b(a[870]), .out(
        \prgm_register/n1742 ) );
  nand2 \prgm_register/C5694  ( .a(\prgm_register/n1741 ), .b(
        \prgm_register/n1742 ), .out(\prgm_register/or_signal [870]) );
  nand2 \prgm_register/C5695  ( .a(enable), .b(a[870]), .out(
        \prgm_register/n1743 ) );
  nand2 \prgm_register/C5696  ( .a(\prgm_register/en_not ), .b(a[871]), .out(
        \prgm_register/n1744 ) );
  nand2 \prgm_register/C5697  ( .a(\prgm_register/n1743 ), .b(
        \prgm_register/n1744 ), .out(\prgm_register/or_signal [871]) );
  nand2 \prgm_register/C5698  ( .a(enable), .b(a[871]), .out(
        \prgm_register/n1745 ) );
  nand2 \prgm_register/C5699  ( .a(\prgm_register/en_not ), .b(a[872]), .out(
        \prgm_register/n1746 ) );
  nand2 \prgm_register/C5700  ( .a(\prgm_register/n1745 ), .b(
        \prgm_register/n1746 ), .out(\prgm_register/or_signal [872]) );
  nand2 \prgm_register/C5701  ( .a(enable), .b(a[872]), .out(
        \prgm_register/n1747 ) );
  nand2 \prgm_register/C5702  ( .a(\prgm_register/en_not ), .b(a[873]), .out(
        \prgm_register/n1748 ) );
  nand2 \prgm_register/C5703  ( .a(\prgm_register/n1747 ), .b(
        \prgm_register/n1748 ), .out(\prgm_register/or_signal [873]) );
  nand2 \prgm_register/C5704  ( .a(enable), .b(a[873]), .out(
        \prgm_register/n1749 ) );
  nand2 \prgm_register/C5705  ( .a(\prgm_register/en_not ), .b(a[874]), .out(
        \prgm_register/n1750 ) );
  nand2 \prgm_register/C5706  ( .a(\prgm_register/n1749 ), .b(
        \prgm_register/n1750 ), .out(\prgm_register/or_signal [874]) );
  nand2 \prgm_register/C5707  ( .a(enable), .b(a[874]), .out(
        \prgm_register/n1751 ) );
  nand2 \prgm_register/C5708  ( .a(\prgm_register/en_not ), .b(a[875]), .out(
        \prgm_register/n1752 ) );
  nand2 \prgm_register/C5709  ( .a(\prgm_register/n1751 ), .b(
        \prgm_register/n1752 ), .out(\prgm_register/or_signal [875]) );
  nand2 \prgm_register/C5710  ( .a(enable), .b(a[875]), .out(
        \prgm_register/n1753 ) );
  nand2 \prgm_register/C5711  ( .a(\prgm_register/en_not ), .b(a[876]), .out(
        \prgm_register/n1754 ) );
  nand2 \prgm_register/C5712  ( .a(\prgm_register/n1753 ), .b(
        \prgm_register/n1754 ), .out(\prgm_register/or_signal [876]) );
  nand2 \prgm_register/C5713  ( .a(enable), .b(a[876]), .out(
        \prgm_register/n1755 ) );
  nand2 \prgm_register/C5714  ( .a(\prgm_register/en_not ), .b(a[877]), .out(
        \prgm_register/n1756 ) );
  nand2 \prgm_register/C5715  ( .a(\prgm_register/n1755 ), .b(
        \prgm_register/n1756 ), .out(\prgm_register/or_signal [877]) );
  nand2 \prgm_register/C5716  ( .a(enable), .b(a[877]), .out(
        \prgm_register/n1757 ) );
  nand2 \prgm_register/C5717  ( .a(\prgm_register/en_not ), .b(a[878]), .out(
        \prgm_register/n1758 ) );
  nand2 \prgm_register/C5718  ( .a(\prgm_register/n1757 ), .b(
        \prgm_register/n1758 ), .out(\prgm_register/or_signal [878]) );
  nand2 \prgm_register/C5719  ( .a(enable), .b(a[878]), .out(
        \prgm_register/n1759 ) );
  nand2 \prgm_register/C5720  ( .a(\prgm_register/en_not ), .b(a[879]), .out(
        \prgm_register/n1760 ) );
  nand2 \prgm_register/C5721  ( .a(\prgm_register/n1759 ), .b(
        \prgm_register/n1760 ), .out(\prgm_register/or_signal [879]) );
  nand2 \prgm_register/C5722  ( .a(enable), .b(a[879]), .out(
        \prgm_register/n1761 ) );
  nand2 \prgm_register/C5723  ( .a(\prgm_register/en_not ), .b(a[880]), .out(
        \prgm_register/n1762 ) );
  nand2 \prgm_register/C5724  ( .a(\prgm_register/n1761 ), .b(
        \prgm_register/n1762 ), .out(\prgm_register/or_signal [880]) );
  nand2 \prgm_register/C5725  ( .a(enable), .b(a[880]), .out(
        \prgm_register/n1763 ) );
  nand2 \prgm_register/C5726  ( .a(\prgm_register/en_not ), .b(a[881]), .out(
        \prgm_register/n1764 ) );
  nand2 \prgm_register/C5727  ( .a(\prgm_register/n1763 ), .b(
        \prgm_register/n1764 ), .out(\prgm_register/or_signal [881]) );
  nand2 \prgm_register/C5728  ( .a(enable), .b(a[881]), .out(
        \prgm_register/n1765 ) );
  nand2 \prgm_register/C5729  ( .a(\prgm_register/en_not ), .b(a[882]), .out(
        \prgm_register/n1766 ) );
  nand2 \prgm_register/C5730  ( .a(\prgm_register/n1765 ), .b(
        \prgm_register/n1766 ), .out(\prgm_register/or_signal [882]) );
  nand2 \prgm_register/C5731  ( .a(enable), .b(a[882]), .out(
        \prgm_register/n1767 ) );
  nand2 \prgm_register/C5732  ( .a(\prgm_register/en_not ), .b(a[883]), .out(
        \prgm_register/n1768 ) );
  nand2 \prgm_register/C5733  ( .a(\prgm_register/n1767 ), .b(
        \prgm_register/n1768 ), .out(\prgm_register/or_signal [883]) );
  nand2 \prgm_register/C5734  ( .a(enable), .b(a[883]), .out(
        \prgm_register/n1769 ) );
  nand2 \prgm_register/C5735  ( .a(\prgm_register/en_not ), .b(a[884]), .out(
        \prgm_register/n1770 ) );
  nand2 \prgm_register/C5736  ( .a(\prgm_register/n1769 ), .b(
        \prgm_register/n1770 ), .out(\prgm_register/or_signal [884]) );
  nand2 \prgm_register/C5737  ( .a(enable), .b(a[884]), .out(
        \prgm_register/n1771 ) );
  nand2 \prgm_register/C5738  ( .a(\prgm_register/en_not ), .b(a[885]), .out(
        \prgm_register/n1772 ) );
  nand2 \prgm_register/C5739  ( .a(\prgm_register/n1771 ), .b(
        \prgm_register/n1772 ), .out(\prgm_register/or_signal [885]) );
  nand2 \prgm_register/C5740  ( .a(enable), .b(a[885]), .out(
        \prgm_register/n1773 ) );
  nand2 \prgm_register/C5741  ( .a(\prgm_register/en_not ), .b(a[886]), .out(
        \prgm_register/n1774 ) );
  nand2 \prgm_register/C5742  ( .a(\prgm_register/n1773 ), .b(
        \prgm_register/n1774 ), .out(\prgm_register/or_signal [886]) );
  nand2 \prgm_register/C5743  ( .a(enable), .b(a[886]), .out(
        \prgm_register/n1775 ) );
  nand2 \prgm_register/C5744  ( .a(\prgm_register/en_not ), .b(a[887]), .out(
        \prgm_register/n1776 ) );
  nand2 \prgm_register/C5745  ( .a(\prgm_register/n1775 ), .b(
        \prgm_register/n1776 ), .out(\prgm_register/or_signal [887]) );
  nand2 \prgm_register/C5746  ( .a(enable), .b(a[887]), .out(
        \prgm_register/n1777 ) );
  nand2 \prgm_register/C5747  ( .a(\prgm_register/en_not ), .b(a[888]), .out(
        \prgm_register/n1778 ) );
  nand2 \prgm_register/C5748  ( .a(\prgm_register/n1777 ), .b(
        \prgm_register/n1778 ), .out(\prgm_register/or_signal [888]) );
  nand2 \prgm_register/C5749  ( .a(enable), .b(a[888]), .out(
        \prgm_register/n1779 ) );
  nand2 \prgm_register/C5750  ( .a(\prgm_register/en_not ), .b(a[889]), .out(
        \prgm_register/n1780 ) );
  nand2 \prgm_register/C5751  ( .a(\prgm_register/n1779 ), .b(
        \prgm_register/n1780 ), .out(\prgm_register/or_signal [889]) );
  nand2 \prgm_register/C5752  ( .a(enable), .b(a[889]), .out(
        \prgm_register/n1781 ) );
  nand2 \prgm_register/C5753  ( .a(\prgm_register/en_not ), .b(a[890]), .out(
        \prgm_register/n1782 ) );
  nand2 \prgm_register/C5754  ( .a(\prgm_register/n1781 ), .b(
        \prgm_register/n1782 ), .out(\prgm_register/or_signal [890]) );
  nand2 \prgm_register/C5755  ( .a(enable), .b(a[890]), .out(
        \prgm_register/n1783 ) );
  nand2 \prgm_register/C5756  ( .a(\prgm_register/en_not ), .b(a[891]), .out(
        \prgm_register/n1784 ) );
  nand2 \prgm_register/C5757  ( .a(\prgm_register/n1783 ), .b(
        \prgm_register/n1784 ), .out(\prgm_register/or_signal [891]) );
  nand2 \prgm_register/C5758  ( .a(enable), .b(a[891]), .out(
        \prgm_register/n1785 ) );
  nand2 \prgm_register/C5759  ( .a(\prgm_register/en_not ), .b(a[892]), .out(
        \prgm_register/n1786 ) );
  nand2 \prgm_register/C5760  ( .a(\prgm_register/n1785 ), .b(
        \prgm_register/n1786 ), .out(\prgm_register/or_signal [892]) );
  nand2 \prgm_register/C5761  ( .a(enable), .b(a[892]), .out(
        \prgm_register/n1787 ) );
  nand2 \prgm_register/C5762  ( .a(\prgm_register/en_not ), .b(a[893]), .out(
        \prgm_register/n1788 ) );
  nand2 \prgm_register/C5763  ( .a(\prgm_register/n1787 ), .b(
        \prgm_register/n1788 ), .out(\prgm_register/or_signal [893]) );
  nand2 \prgm_register/C5764  ( .a(enable), .b(a[893]), .out(
        \prgm_register/n1789 ) );
  nand2 \prgm_register/C5765  ( .a(\prgm_register/en_not ), .b(a[894]), .out(
        \prgm_register/n1790 ) );
  nand2 \prgm_register/C5766  ( .a(\prgm_register/n1789 ), .b(
        \prgm_register/n1790 ), .out(\prgm_register/or_signal [894]) );
  nand2 \prgm_register/C5767  ( .a(enable), .b(a[894]), .out(
        \prgm_register/n1791 ) );
  nand2 \prgm_register/C5768  ( .a(\prgm_register/en_not ), .b(a[895]), .out(
        \prgm_register/n1792 ) );
  nand2 \prgm_register/C5769  ( .a(\prgm_register/n1791 ), .b(
        \prgm_register/n1792 ), .out(\prgm_register/or_signal [895]) );
  nand2 \prgm_register/C5770  ( .a(enable), .b(a[895]), .out(
        \prgm_register/n1793 ) );
  nand2 \prgm_register/C5771  ( .a(\prgm_register/en_not ), .b(a[896]), .out(
        \prgm_register/n1794 ) );
  nand2 \prgm_register/C5772  ( .a(\prgm_register/n1793 ), .b(
        \prgm_register/n1794 ), .out(\prgm_register/or_signal [896]) );
  nand2 \prgm_register/C5773  ( .a(enable), .b(a[896]), .out(
        \prgm_register/n1795 ) );
  nand2 \prgm_register/C5774  ( .a(\prgm_register/en_not ), .b(a[897]), .out(
        \prgm_register/n1796 ) );
  nand2 \prgm_register/C5775  ( .a(\prgm_register/n1795 ), .b(
        \prgm_register/n1796 ), .out(\prgm_register/or_signal [897]) );
  nand2 \prgm_register/C5776  ( .a(enable), .b(a[897]), .out(
        \prgm_register/n1797 ) );
  nand2 \prgm_register/C5777  ( .a(\prgm_register/en_not ), .b(a[898]), .out(
        \prgm_register/n1798 ) );
  nand2 \prgm_register/C5778  ( .a(\prgm_register/n1797 ), .b(
        \prgm_register/n1798 ), .out(\prgm_register/or_signal [898]) );
  nand2 \prgm_register/C5779  ( .a(enable), .b(a[898]), .out(
        \prgm_register/n1799 ) );
  nand2 \prgm_register/C5780  ( .a(\prgm_register/en_not ), .b(a[899]), .out(
        \prgm_register/n1800 ) );
  nand2 \prgm_register/C5781  ( .a(\prgm_register/n1799 ), .b(
        \prgm_register/n1800 ), .out(\prgm_register/or_signal [899]) );
  nand2 \prgm_register/C5782  ( .a(enable), .b(a[899]), .out(
        \prgm_register/n1801 ) );
  nand2 \prgm_register/C5783  ( .a(\prgm_register/en_not ), .b(a[900]), .out(
        \prgm_register/n1802 ) );
  nand2 \prgm_register/C5784  ( .a(\prgm_register/n1801 ), .b(
        \prgm_register/n1802 ), .out(\prgm_register/or_signal [900]) );
  nand2 \prgm_register/C5785  ( .a(enable), .b(a[900]), .out(
        \prgm_register/n1803 ) );
  nand2 \prgm_register/C5786  ( .a(\prgm_register/en_not ), .b(a[901]), .out(
        \prgm_register/n1804 ) );
  nand2 \prgm_register/C5787  ( .a(\prgm_register/n1803 ), .b(
        \prgm_register/n1804 ), .out(\prgm_register/or_signal [901]) );
  nand2 \prgm_register/C5788  ( .a(enable), .b(a[901]), .out(
        \prgm_register/n1805 ) );
  nand2 \prgm_register/C5789  ( .a(\prgm_register/en_not ), .b(a[902]), .out(
        \prgm_register/n1806 ) );
  nand2 \prgm_register/C5790  ( .a(\prgm_register/n1805 ), .b(
        \prgm_register/n1806 ), .out(\prgm_register/or_signal [902]) );
  nand2 \prgm_register/C5791  ( .a(enable), .b(a[902]), .out(
        \prgm_register/n1807 ) );
  nand2 \prgm_register/C5792  ( .a(\prgm_register/en_not ), .b(a[903]), .out(
        \prgm_register/n1808 ) );
  nand2 \prgm_register/C5793  ( .a(\prgm_register/n1807 ), .b(
        \prgm_register/n1808 ), .out(\prgm_register/or_signal [903]) );
  nand2 \prgm_register/C5794  ( .a(enable), .b(a[903]), .out(
        \prgm_register/n1809 ) );
  nand2 \prgm_register/C5795  ( .a(\prgm_register/en_not ), .b(a[904]), .out(
        \prgm_register/n1810 ) );
  nand2 \prgm_register/C5796  ( .a(\prgm_register/n1809 ), .b(
        \prgm_register/n1810 ), .out(\prgm_register/or_signal [904]) );
  nand2 \prgm_register/C5797  ( .a(enable), .b(a[904]), .out(
        \prgm_register/n1811 ) );
  nand2 \prgm_register/C5798  ( .a(\prgm_register/en_not ), .b(a[905]), .out(
        \prgm_register/n1812 ) );
  nand2 \prgm_register/C5799  ( .a(\prgm_register/n1811 ), .b(
        \prgm_register/n1812 ), .out(\prgm_register/or_signal [905]) );
  nand2 \prgm_register/C5800  ( .a(enable), .b(a[905]), .out(
        \prgm_register/n1813 ) );
  nand2 \prgm_register/C5801  ( .a(\prgm_register/en_not ), .b(a[906]), .out(
        \prgm_register/n1814 ) );
  nand2 \prgm_register/C5802  ( .a(\prgm_register/n1813 ), .b(
        \prgm_register/n1814 ), .out(\prgm_register/or_signal [906]) );
  nand2 \prgm_register/C5803  ( .a(enable), .b(a[906]), .out(
        \prgm_register/n1815 ) );
  nand2 \prgm_register/C5804  ( .a(\prgm_register/en_not ), .b(a[907]), .out(
        \prgm_register/n1816 ) );
  nand2 \prgm_register/C5805  ( .a(\prgm_register/n1815 ), .b(
        \prgm_register/n1816 ), .out(\prgm_register/or_signal [907]) );
  nand2 \prgm_register/C5806  ( .a(enable), .b(a[907]), .out(
        \prgm_register/n1817 ) );
  nand2 \prgm_register/C5807  ( .a(\prgm_register/en_not ), .b(a[908]), .out(
        \prgm_register/n1818 ) );
  nand2 \prgm_register/C5808  ( .a(\prgm_register/n1817 ), .b(
        \prgm_register/n1818 ), .out(\prgm_register/or_signal [908]) );
  nand2 \prgm_register/C5809  ( .a(enable), .b(a[908]), .out(
        \prgm_register/n1819 ) );
  nand2 \prgm_register/C5810  ( .a(\prgm_register/en_not ), .b(a[909]), .out(
        \prgm_register/n1820 ) );
  nand2 \prgm_register/C5811  ( .a(\prgm_register/n1819 ), .b(
        \prgm_register/n1820 ), .out(\prgm_register/or_signal [909]) );
  nand2 \prgm_register/C5812  ( .a(enable), .b(a[909]), .out(
        \prgm_register/n1821 ) );
  nand2 \prgm_register/C5813  ( .a(\prgm_register/en_not ), .b(a[910]), .out(
        \prgm_register/n1822 ) );
  nand2 \prgm_register/C5814  ( .a(\prgm_register/n1821 ), .b(
        \prgm_register/n1822 ), .out(\prgm_register/or_signal [910]) );
  nand2 \prgm_register/C5815  ( .a(enable), .b(a[910]), .out(
        \prgm_register/n1823 ) );
  nand2 \prgm_register/C5816  ( .a(\prgm_register/en_not ), .b(a[911]), .out(
        \prgm_register/n1824 ) );
  nand2 \prgm_register/C5817  ( .a(\prgm_register/n1823 ), .b(
        \prgm_register/n1824 ), .out(\prgm_register/or_signal [911]) );
  nand2 \prgm_register/C5818  ( .a(enable), .b(a[911]), .out(
        \prgm_register/n1825 ) );
  nand2 \prgm_register/C5819  ( .a(\prgm_register/en_not ), .b(a[912]), .out(
        \prgm_register/n1826 ) );
  nand2 \prgm_register/C5820  ( .a(\prgm_register/n1825 ), .b(
        \prgm_register/n1826 ), .out(\prgm_register/or_signal [912]) );
  nand2 \prgm_register/C5821  ( .a(enable), .b(a[912]), .out(
        \prgm_register/n1827 ) );
  nand2 \prgm_register/C5822  ( .a(\prgm_register/en_not ), .b(a[913]), .out(
        \prgm_register/n1828 ) );
  nand2 \prgm_register/C5823  ( .a(\prgm_register/n1827 ), .b(
        \prgm_register/n1828 ), .out(\prgm_register/or_signal [913]) );
  nand2 \prgm_register/C5824  ( .a(enable), .b(a[913]), .out(
        \prgm_register/n1829 ) );
  nand2 \prgm_register/C5825  ( .a(\prgm_register/en_not ), .b(a[914]), .out(
        \prgm_register/n1830 ) );
  nand2 \prgm_register/C5826  ( .a(\prgm_register/n1829 ), .b(
        \prgm_register/n1830 ), .out(\prgm_register/or_signal [914]) );
  nand2 \prgm_register/C5827  ( .a(enable), .b(a[914]), .out(
        \prgm_register/n1831 ) );
  nand2 \prgm_register/C5828  ( .a(\prgm_register/en_not ), .b(a[915]), .out(
        \prgm_register/n1832 ) );
  nand2 \prgm_register/C5829  ( .a(\prgm_register/n1831 ), .b(
        \prgm_register/n1832 ), .out(\prgm_register/or_signal [915]) );
  nand2 \prgm_register/C5830  ( .a(enable), .b(a[915]), .out(
        \prgm_register/n1833 ) );
  nand2 \prgm_register/C5831  ( .a(\prgm_register/en_not ), .b(a[916]), .out(
        \prgm_register/n1834 ) );
  nand2 \prgm_register/C5832  ( .a(\prgm_register/n1833 ), .b(
        \prgm_register/n1834 ), .out(\prgm_register/or_signal [916]) );
  nand2 \prgm_register/C5833  ( .a(enable), .b(a[916]), .out(
        \prgm_register/n1835 ) );
  nand2 \prgm_register/C5834  ( .a(\prgm_register/en_not ), .b(a[917]), .out(
        \prgm_register/n1836 ) );
  nand2 \prgm_register/C5835  ( .a(\prgm_register/n1835 ), .b(
        \prgm_register/n1836 ), .out(\prgm_register/or_signal [917]) );
  nand2 \prgm_register/C5836  ( .a(enable), .b(a[917]), .out(
        \prgm_register/n1837 ) );
  nand2 \prgm_register/C5837  ( .a(\prgm_register/en_not ), .b(a[918]), .out(
        \prgm_register/n1838 ) );
  nand2 \prgm_register/C5838  ( .a(\prgm_register/n1837 ), .b(
        \prgm_register/n1838 ), .out(\prgm_register/or_signal [918]) );
  nand2 \prgm_register/C5839  ( .a(enable), .b(a[918]), .out(
        \prgm_register/n1839 ) );
  nand2 \prgm_register/C5840  ( .a(\prgm_register/en_not ), .b(a[919]), .out(
        \prgm_register/n1840 ) );
  nand2 \prgm_register/C5841  ( .a(\prgm_register/n1839 ), .b(
        \prgm_register/n1840 ), .out(\prgm_register/or_signal [919]) );
  nand2 \prgm_register/C5842  ( .a(enable), .b(a[919]), .out(
        \prgm_register/n1841 ) );
  nand2 \prgm_register/C5843  ( .a(\prgm_register/en_not ), .b(a[920]), .out(
        \prgm_register/n1842 ) );
  nand2 \prgm_register/C5844  ( .a(\prgm_register/n1841 ), .b(
        \prgm_register/n1842 ), .out(\prgm_register/or_signal [920]) );
  nand2 \prgm_register/C5845  ( .a(enable), .b(a[920]), .out(
        \prgm_register/n1843 ) );
  nand2 \prgm_register/C5846  ( .a(\prgm_register/en_not ), .b(a[921]), .out(
        \prgm_register/n1844 ) );
  nand2 \prgm_register/C5847  ( .a(\prgm_register/n1843 ), .b(
        \prgm_register/n1844 ), .out(\prgm_register/or_signal [921]) );
  nand2 \prgm_register/C5848  ( .a(enable), .b(a[921]), .out(
        \prgm_register/n1845 ) );
  nand2 \prgm_register/C5849  ( .a(\prgm_register/en_not ), .b(a[922]), .out(
        \prgm_register/n1846 ) );
  nand2 \prgm_register/C5850  ( .a(\prgm_register/n1845 ), .b(
        \prgm_register/n1846 ), .out(\prgm_register/or_signal [922]) );
  nand2 \prgm_register/C5851  ( .a(enable), .b(a[922]), .out(
        \prgm_register/n1847 ) );
  nand2 \prgm_register/C5852  ( .a(\prgm_register/en_not ), .b(a[923]), .out(
        \prgm_register/n1848 ) );
  nand2 \prgm_register/C5853  ( .a(\prgm_register/n1847 ), .b(
        \prgm_register/n1848 ), .out(\prgm_register/or_signal [923]) );
  nand2 \prgm_register/C5854  ( .a(enable), .b(a[923]), .out(
        \prgm_register/n1849 ) );
  nand2 \prgm_register/C5855  ( .a(\prgm_register/en_not ), .b(a[924]), .out(
        \prgm_register/n1850 ) );
  nand2 \prgm_register/C5856  ( .a(\prgm_register/n1849 ), .b(
        \prgm_register/n1850 ), .out(\prgm_register/or_signal [924]) );
  nand2 \prgm_register/C5857  ( .a(enable), .b(a[924]), .out(
        \prgm_register/n1851 ) );
  nand2 \prgm_register/C5858  ( .a(\prgm_register/en_not ), .b(a[925]), .out(
        \prgm_register/n1852 ) );
  nand2 \prgm_register/C5859  ( .a(\prgm_register/n1851 ), .b(
        \prgm_register/n1852 ), .out(\prgm_register/or_signal [925]) );
  nand2 \prgm_register/C5860  ( .a(enable), .b(a[925]), .out(
        \prgm_register/n1853 ) );
  nand2 \prgm_register/C5861  ( .a(\prgm_register/en_not ), .b(a[926]), .out(
        \prgm_register/n1854 ) );
  nand2 \prgm_register/C5862  ( .a(\prgm_register/n1853 ), .b(
        \prgm_register/n1854 ), .out(\prgm_register/or_signal [926]) );
  nand2 \prgm_register/C5863  ( .a(enable), .b(a[926]), .out(
        \prgm_register/n1855 ) );
  nand2 \prgm_register/C5864  ( .a(\prgm_register/en_not ), .b(a[927]), .out(
        \prgm_register/n1856 ) );
  nand2 \prgm_register/C5865  ( .a(\prgm_register/n1855 ), .b(
        \prgm_register/n1856 ), .out(\prgm_register/or_signal [927]) );
  nand2 \prgm_register/C5866  ( .a(enable), .b(a[927]), .out(
        \prgm_register/n1857 ) );
  nand2 \prgm_register/C5867  ( .a(\prgm_register/en_not ), .b(a[928]), .out(
        \prgm_register/n1858 ) );
  nand2 \prgm_register/C5868  ( .a(\prgm_register/n1857 ), .b(
        \prgm_register/n1858 ), .out(\prgm_register/or_signal [928]) );
  nand2 \prgm_register/C5869  ( .a(enable), .b(a[928]), .out(
        \prgm_register/n1859 ) );
  nand2 \prgm_register/C5870  ( .a(\prgm_register/en_not ), .b(a[929]), .out(
        \prgm_register/n1860 ) );
  nand2 \prgm_register/C5871  ( .a(\prgm_register/n1859 ), .b(
        \prgm_register/n1860 ), .out(\prgm_register/or_signal [929]) );
  nand2 \prgm_register/C5872  ( .a(enable), .b(a[929]), .out(
        \prgm_register/n1861 ) );
  nand2 \prgm_register/C5873  ( .a(\prgm_register/en_not ), .b(a[930]), .out(
        \prgm_register/n1862 ) );
  nand2 \prgm_register/C5874  ( .a(\prgm_register/n1861 ), .b(
        \prgm_register/n1862 ), .out(\prgm_register/or_signal [930]) );
  nand2 \prgm_register/C5875  ( .a(enable), .b(a[930]), .out(
        \prgm_register/n1863 ) );
  nand2 \prgm_register/C5876  ( .a(\prgm_register/en_not ), .b(a[931]), .out(
        \prgm_register/n1864 ) );
  nand2 \prgm_register/C5877  ( .a(\prgm_register/n1863 ), .b(
        \prgm_register/n1864 ), .out(\prgm_register/or_signal [931]) );
  nand2 \prgm_register/C5878  ( .a(enable), .b(a[931]), .out(
        \prgm_register/n1865 ) );
  nand2 \prgm_register/C5879  ( .a(\prgm_register/en_not ), .b(a[932]), .out(
        \prgm_register/n1866 ) );
  nand2 \prgm_register/C5880  ( .a(\prgm_register/n1865 ), .b(
        \prgm_register/n1866 ), .out(\prgm_register/or_signal [932]) );
  nand2 \prgm_register/C5881  ( .a(enable), .b(a[932]), .out(
        \prgm_register/n1867 ) );
  nand2 \prgm_register/C5882  ( .a(\prgm_register/en_not ), .b(a[933]), .out(
        \prgm_register/n1868 ) );
  nand2 \prgm_register/C5883  ( .a(\prgm_register/n1867 ), .b(
        \prgm_register/n1868 ), .out(\prgm_register/or_signal [933]) );
  nand2 \prgm_register/C5884  ( .a(enable), .b(a[933]), .out(
        \prgm_register/n1869 ) );
  nand2 \prgm_register/C5885  ( .a(\prgm_register/en_not ), .b(a[934]), .out(
        \prgm_register/n1870 ) );
  nand2 \prgm_register/C5886  ( .a(\prgm_register/n1869 ), .b(
        \prgm_register/n1870 ), .out(\prgm_register/or_signal [934]) );
  nand2 \prgm_register/C5887  ( .a(enable), .b(a[934]), .out(
        \prgm_register/n1871 ) );
  nand2 \prgm_register/C5888  ( .a(\prgm_register/en_not ), .b(a[935]), .out(
        \prgm_register/n1872 ) );
  nand2 \prgm_register/C5889  ( .a(\prgm_register/n1871 ), .b(
        \prgm_register/n1872 ), .out(\prgm_register/or_signal [935]) );
  nand2 \prgm_register/C5890  ( .a(enable), .b(a[935]), .out(
        \prgm_register/n1873 ) );
  nand2 \prgm_register/C5891  ( .a(\prgm_register/en_not ), .b(a[936]), .out(
        \prgm_register/n1874 ) );
  nand2 \prgm_register/C5892  ( .a(\prgm_register/n1873 ), .b(
        \prgm_register/n1874 ), .out(\prgm_register/or_signal [936]) );
  nand2 \prgm_register/C5893  ( .a(enable), .b(a[936]), .out(
        \prgm_register/n1875 ) );
  nand2 \prgm_register/C5894  ( .a(\prgm_register/en_not ), .b(a[937]), .out(
        \prgm_register/n1876 ) );
  nand2 \prgm_register/C5895  ( .a(\prgm_register/n1875 ), .b(
        \prgm_register/n1876 ), .out(\prgm_register/or_signal [937]) );
  nand2 \prgm_register/C5896  ( .a(enable), .b(a[937]), .out(
        \prgm_register/n1877 ) );
  nand2 \prgm_register/C5897  ( .a(\prgm_register/en_not ), .b(a[938]), .out(
        \prgm_register/n1878 ) );
  nand2 \prgm_register/C5898  ( .a(\prgm_register/n1877 ), .b(
        \prgm_register/n1878 ), .out(\prgm_register/or_signal [938]) );
  nand2 \prgm_register/C5899  ( .a(enable), .b(a[938]), .out(
        \prgm_register/n1879 ) );
  nand2 \prgm_register/C5900  ( .a(\prgm_register/en_not ), .b(a[939]), .out(
        \prgm_register/n1880 ) );
  nand2 \prgm_register/C5901  ( .a(\prgm_register/n1879 ), .b(
        \prgm_register/n1880 ), .out(\prgm_register/or_signal [939]) );
  nand2 \prgm_register/C5902  ( .a(enable), .b(a[939]), .out(
        \prgm_register/n1881 ) );
  nand2 \prgm_register/C5903  ( .a(\prgm_register/en_not ), .b(a[940]), .out(
        \prgm_register/n1882 ) );
  nand2 \prgm_register/C5904  ( .a(\prgm_register/n1881 ), .b(
        \prgm_register/n1882 ), .out(\prgm_register/or_signal [940]) );
  nand2 \prgm_register/C5905  ( .a(enable), .b(a[940]), .out(
        \prgm_register/n1883 ) );
  nand2 \prgm_register/C5906  ( .a(\prgm_register/en_not ), .b(a[941]), .out(
        \prgm_register/n1884 ) );
  nand2 \prgm_register/C5907  ( .a(\prgm_register/n1883 ), .b(
        \prgm_register/n1884 ), .out(\prgm_register/or_signal [941]) );
  nand2 \prgm_register/C5908  ( .a(enable), .b(a[941]), .out(
        \prgm_register/n1885 ) );
  nand2 \prgm_register/C5909  ( .a(\prgm_register/en_not ), .b(a[942]), .out(
        \prgm_register/n1886 ) );
  nand2 \prgm_register/C5910  ( .a(\prgm_register/n1885 ), .b(
        \prgm_register/n1886 ), .out(\prgm_register/or_signal [942]) );
  nand2 \prgm_register/C5911  ( .a(enable), .b(a[942]), .out(
        \prgm_register/n1887 ) );
  nand2 \prgm_register/C5912  ( .a(\prgm_register/en_not ), .b(a[943]), .out(
        \prgm_register/n1888 ) );
  nand2 \prgm_register/C5913  ( .a(\prgm_register/n1887 ), .b(
        \prgm_register/n1888 ), .out(\prgm_register/or_signal [943]) );
  nand2 \prgm_register/C5914  ( .a(enable), .b(a[943]), .out(
        \prgm_register/n1889 ) );
  nand2 \prgm_register/C5915  ( .a(\prgm_register/en_not ), .b(a[944]), .out(
        \prgm_register/n1890 ) );
  nand2 \prgm_register/C5916  ( .a(\prgm_register/n1889 ), .b(
        \prgm_register/n1890 ), .out(\prgm_register/or_signal [944]) );
  nand2 \prgm_register/C5917  ( .a(enable), .b(a[944]), .out(
        \prgm_register/n1891 ) );
  nand2 \prgm_register/C5918  ( .a(\prgm_register/en_not ), .b(a[945]), .out(
        \prgm_register/n1892 ) );
  nand2 \prgm_register/C5919  ( .a(\prgm_register/n1891 ), .b(
        \prgm_register/n1892 ), .out(\prgm_register/or_signal [945]) );
  nand2 \prgm_register/C5920  ( .a(enable), .b(a[945]), .out(
        \prgm_register/n1893 ) );
  nand2 \prgm_register/C5921  ( .a(\prgm_register/en_not ), .b(a[946]), .out(
        \prgm_register/n1894 ) );
  nand2 \prgm_register/C5922  ( .a(\prgm_register/n1893 ), .b(
        \prgm_register/n1894 ), .out(\prgm_register/or_signal [946]) );
  nand2 \prgm_register/C5923  ( .a(enable), .b(a[946]), .out(
        \prgm_register/n1895 ) );
  nand2 \prgm_register/C5924  ( .a(\prgm_register/en_not ), .b(a[947]), .out(
        \prgm_register/n1896 ) );
  nand2 \prgm_register/C5925  ( .a(\prgm_register/n1895 ), .b(
        \prgm_register/n1896 ), .out(\prgm_register/or_signal [947]) );
  nand2 \prgm_register/C5926  ( .a(enable), .b(a[947]), .out(
        \prgm_register/n1897 ) );
  nand2 \prgm_register/C5927  ( .a(\prgm_register/en_not ), .b(a[948]), .out(
        \prgm_register/n1898 ) );
  nand2 \prgm_register/C5928  ( .a(\prgm_register/n1897 ), .b(
        \prgm_register/n1898 ), .out(\prgm_register/or_signal [948]) );
  nand2 \prgm_register/C5929  ( .a(enable), .b(a[948]), .out(
        \prgm_register/n1899 ) );
  nand2 \prgm_register/C5930  ( .a(\prgm_register/en_not ), .b(a[949]), .out(
        \prgm_register/n1900 ) );
  nand2 \prgm_register/C5931  ( .a(\prgm_register/n1899 ), .b(
        \prgm_register/n1900 ), .out(\prgm_register/or_signal [949]) );
  nand2 \prgm_register/C5932  ( .a(enable), .b(a[949]), .out(
        \prgm_register/n1901 ) );
  nand2 \prgm_register/C5933  ( .a(\prgm_register/en_not ), .b(a[950]), .out(
        \prgm_register/n1902 ) );
  nand2 \prgm_register/C5934  ( .a(\prgm_register/n1901 ), .b(
        \prgm_register/n1902 ), .out(\prgm_register/or_signal [950]) );
  nand2 \prgm_register/C5935  ( .a(enable), .b(a[950]), .out(
        \prgm_register/n1903 ) );
  nand2 \prgm_register/C5936  ( .a(\prgm_register/en_not ), .b(a[951]), .out(
        \prgm_register/n1904 ) );
  nand2 \prgm_register/C5937  ( .a(\prgm_register/n1903 ), .b(
        \prgm_register/n1904 ), .out(\prgm_register/or_signal [951]) );
  nand2 \prgm_register/C5938  ( .a(enable), .b(a[951]), .out(
        \prgm_register/n1905 ) );
  nand2 \prgm_register/C5939  ( .a(\prgm_register/en_not ), .b(a[952]), .out(
        \prgm_register/n1906 ) );
  nand2 \prgm_register/C5940  ( .a(\prgm_register/n1905 ), .b(
        \prgm_register/n1906 ), .out(\prgm_register/or_signal [952]) );
  nand2 \prgm_register/C5941  ( .a(enable), .b(a[952]), .out(
        \prgm_register/n1907 ) );
  nand2 \prgm_register/C5942  ( .a(\prgm_register/en_not ), .b(a[953]), .out(
        \prgm_register/n1908 ) );
  nand2 \prgm_register/C5943  ( .a(\prgm_register/n1907 ), .b(
        \prgm_register/n1908 ), .out(\prgm_register/or_signal [953]) );
  nand2 \prgm_register/C5944  ( .a(enable), .b(a[953]), .out(
        \prgm_register/n1909 ) );
  nand2 \prgm_register/C5945  ( .a(\prgm_register/en_not ), .b(a[954]), .out(
        \prgm_register/n1910 ) );
  nand2 \prgm_register/C5946  ( .a(\prgm_register/n1909 ), .b(
        \prgm_register/n1910 ), .out(\prgm_register/or_signal [954]) );
  nand2 \prgm_register/C5947  ( .a(enable), .b(a[954]), .out(
        \prgm_register/n1911 ) );
  nand2 \prgm_register/C5948  ( .a(\prgm_register/en_not ), .b(a[955]), .out(
        \prgm_register/n1912 ) );
  nand2 \prgm_register/C5949  ( .a(\prgm_register/n1911 ), .b(
        \prgm_register/n1912 ), .out(\prgm_register/or_signal [955]) );
  nand2 \prgm_register/C5950  ( .a(enable), .b(a[955]), .out(
        \prgm_register/n1913 ) );
  nand2 \prgm_register/C5951  ( .a(\prgm_register/en_not ), .b(a[956]), .out(
        \prgm_register/n1914 ) );
  nand2 \prgm_register/C5952  ( .a(\prgm_register/n1913 ), .b(
        \prgm_register/n1914 ), .out(\prgm_register/or_signal [956]) );
  nand2 \prgm_register/C5953  ( .a(enable), .b(a[956]), .out(
        \prgm_register/n1915 ) );
  nand2 \prgm_register/C5954  ( .a(\prgm_register/en_not ), .b(a[957]), .out(
        \prgm_register/n1916 ) );
  nand2 \prgm_register/C5955  ( .a(\prgm_register/n1915 ), .b(
        \prgm_register/n1916 ), .out(\prgm_register/or_signal [957]) );
  nand2 \prgm_register/C5956  ( .a(enable), .b(a[957]), .out(
        \prgm_register/n1917 ) );
  nand2 \prgm_register/C5957  ( .a(\prgm_register/en_not ), .b(a[958]), .out(
        \prgm_register/n1918 ) );
  nand2 \prgm_register/C5958  ( .a(\prgm_register/n1917 ), .b(
        \prgm_register/n1918 ), .out(\prgm_register/or_signal [958]) );
  nand2 \prgm_register/C5959  ( .a(enable), .b(a[958]), .out(
        \prgm_register/n1919 ) );
  nand2 \prgm_register/C5960  ( .a(\prgm_register/en_not ), .b(a[959]), .out(
        \prgm_register/n1920 ) );
  nand2 \prgm_register/C5961  ( .a(\prgm_register/n1919 ), .b(
        \prgm_register/n1920 ), .out(\prgm_register/or_signal [959]) );
  nand2 \prgm_register/C5962  ( .a(enable), .b(a[959]), .out(
        \prgm_register/n1921 ) );
  nand2 \prgm_register/C5963  ( .a(\prgm_register/en_not ), .b(a[960]), .out(
        \prgm_register/n1922 ) );
  nand2 \prgm_register/C5964  ( .a(\prgm_register/n1921 ), .b(
        \prgm_register/n1922 ), .out(\prgm_register/or_signal [960]) );
  nand2 \prgm_register/C5965  ( .a(enable), .b(a[960]), .out(
        \prgm_register/n1923 ) );
  nand2 \prgm_register/C5966  ( .a(\prgm_register/en_not ), .b(a[961]), .out(
        \prgm_register/n1924 ) );
  nand2 \prgm_register/C5967  ( .a(\prgm_register/n1923 ), .b(
        \prgm_register/n1924 ), .out(\prgm_register/or_signal [961]) );
  nand2 \prgm_register/C5968  ( .a(enable), .b(a[961]), .out(
        \prgm_register/n1925 ) );
  nand2 \prgm_register/C5969  ( .a(\prgm_register/en_not ), .b(a[962]), .out(
        \prgm_register/n1926 ) );
  nand2 \prgm_register/C5970  ( .a(\prgm_register/n1925 ), .b(
        \prgm_register/n1926 ), .out(\prgm_register/or_signal [962]) );
  nand2 \prgm_register/C5971  ( .a(enable), .b(a[962]), .out(
        \prgm_register/n1927 ) );
  nand2 \prgm_register/C5972  ( .a(\prgm_register/en_not ), .b(a[963]), .out(
        \prgm_register/n1928 ) );
  nand2 \prgm_register/C5973  ( .a(\prgm_register/n1927 ), .b(
        \prgm_register/n1928 ), .out(\prgm_register/or_signal [963]) );
  nand2 \prgm_register/C5974  ( .a(enable), .b(a[963]), .out(
        \prgm_register/n1929 ) );
  nand2 \prgm_register/C5975  ( .a(\prgm_register/en_not ), .b(a[964]), .out(
        \prgm_register/n1930 ) );
  nand2 \prgm_register/C5976  ( .a(\prgm_register/n1929 ), .b(
        \prgm_register/n1930 ), .out(\prgm_register/or_signal [964]) );
  nand2 \prgm_register/C5977  ( .a(enable), .b(a[964]), .out(
        \prgm_register/n1931 ) );
  nand2 \prgm_register/C5978  ( .a(\prgm_register/en_not ), .b(a[965]), .out(
        \prgm_register/n1932 ) );
  nand2 \prgm_register/C5979  ( .a(\prgm_register/n1931 ), .b(
        \prgm_register/n1932 ), .out(\prgm_register/or_signal [965]) );
  nand2 \prgm_register/C5980  ( .a(enable), .b(a[965]), .out(
        \prgm_register/n1933 ) );
  nand2 \prgm_register/C5981  ( .a(\prgm_register/en_not ), .b(a[966]), .out(
        \prgm_register/n1934 ) );
  nand2 \prgm_register/C5982  ( .a(\prgm_register/n1933 ), .b(
        \prgm_register/n1934 ), .out(\prgm_register/or_signal [966]) );
  nand2 \prgm_register/C5983  ( .a(enable), .b(a[966]), .out(
        \prgm_register/n1935 ) );
  nand2 \prgm_register/C5984  ( .a(\prgm_register/en_not ), .b(a[967]), .out(
        \prgm_register/n1936 ) );
  nand2 \prgm_register/C5985  ( .a(\prgm_register/n1935 ), .b(
        \prgm_register/n1936 ), .out(\prgm_register/or_signal [967]) );
  nand2 \prgm_register/C5986  ( .a(enable), .b(a[967]), .out(
        \prgm_register/n1937 ) );
  nand2 \prgm_register/C5987  ( .a(\prgm_register/en_not ), .b(a[968]), .out(
        \prgm_register/n1938 ) );
  nand2 \prgm_register/C5988  ( .a(\prgm_register/n1937 ), .b(
        \prgm_register/n1938 ), .out(\prgm_register/or_signal [968]) );
  nand2 \prgm_register/C5989  ( .a(enable), .b(a[968]), .out(
        \prgm_register/n1939 ) );
  nand2 \prgm_register/C5990  ( .a(\prgm_register/en_not ), .b(a[969]), .out(
        \prgm_register/n1940 ) );
  nand2 \prgm_register/C5991  ( .a(\prgm_register/n1939 ), .b(
        \prgm_register/n1940 ), .out(\prgm_register/or_signal [969]) );
  nand2 \prgm_register/C5992  ( .a(enable), .b(a[969]), .out(
        \prgm_register/n1941 ) );
  nand2 \prgm_register/C5993  ( .a(\prgm_register/en_not ), .b(a[970]), .out(
        \prgm_register/n1942 ) );
  nand2 \prgm_register/C5994  ( .a(\prgm_register/n1941 ), .b(
        \prgm_register/n1942 ), .out(\prgm_register/or_signal [970]) );
  nand2 \prgm_register/C5995  ( .a(enable), .b(a[970]), .out(
        \prgm_register/n1943 ) );
  nand2 \prgm_register/C5996  ( .a(\prgm_register/en_not ), .b(a[971]), .out(
        \prgm_register/n1944 ) );
  nand2 \prgm_register/C5997  ( .a(\prgm_register/n1943 ), .b(
        \prgm_register/n1944 ), .out(\prgm_register/or_signal [971]) );
  nand2 \prgm_register/C5998  ( .a(enable), .b(a[971]), .out(
        \prgm_register/n1945 ) );
  nand2 \prgm_register/C5999  ( .a(\prgm_register/en_not ), .b(a[972]), .out(
        \prgm_register/n1946 ) );
  nand2 \prgm_register/C6000  ( .a(\prgm_register/n1945 ), .b(
        \prgm_register/n1946 ), .out(\prgm_register/or_signal [972]) );
  nand2 \prgm_register/C6001  ( .a(enable), .b(a[972]), .out(
        \prgm_register/n1947 ) );
  nand2 \prgm_register/C6002  ( .a(\prgm_register/en_not ), .b(a[973]), .out(
        \prgm_register/n1948 ) );
  nand2 \prgm_register/C6003  ( .a(\prgm_register/n1947 ), .b(
        \prgm_register/n1948 ), .out(\prgm_register/or_signal [973]) );
  nand2 \prgm_register/C6004  ( .a(enable), .b(a[973]), .out(
        \prgm_register/n1949 ) );
  nand2 \prgm_register/C6005  ( .a(\prgm_register/en_not ), .b(a[974]), .out(
        \prgm_register/n1950 ) );
  nand2 \prgm_register/C6006  ( .a(\prgm_register/n1949 ), .b(
        \prgm_register/n1950 ), .out(\prgm_register/or_signal [974]) );
  nand2 \prgm_register/C6007  ( .a(enable), .b(a[974]), .out(
        \prgm_register/n1951 ) );
  nand2 \prgm_register/C6008  ( .a(\prgm_register/en_not ), .b(a[975]), .out(
        \prgm_register/n1952 ) );
  nand2 \prgm_register/C6009  ( .a(\prgm_register/n1951 ), .b(
        \prgm_register/n1952 ), .out(\prgm_register/or_signal [975]) );
  nand2 \prgm_register/C6010  ( .a(enable), .b(a[975]), .out(
        \prgm_register/n1953 ) );
  nand2 \prgm_register/C6011  ( .a(\prgm_register/en_not ), .b(a[976]), .out(
        \prgm_register/n1954 ) );
  nand2 \prgm_register/C6012  ( .a(\prgm_register/n1953 ), .b(
        \prgm_register/n1954 ), .out(\prgm_register/or_signal [976]) );
  nand2 \prgm_register/C6013  ( .a(enable), .b(a[976]), .out(
        \prgm_register/n1955 ) );
  nand2 \prgm_register/C6014  ( .a(\prgm_register/en_not ), .b(a[977]), .out(
        \prgm_register/n1956 ) );
  nand2 \prgm_register/C6015  ( .a(\prgm_register/n1955 ), .b(
        \prgm_register/n1956 ), .out(\prgm_register/or_signal [977]) );
  nand2 \prgm_register/C6016  ( .a(enable), .b(a[977]), .out(
        \prgm_register/n1957 ) );
  nand2 \prgm_register/C6017  ( .a(\prgm_register/en_not ), .b(a[978]), .out(
        \prgm_register/n1958 ) );
  nand2 \prgm_register/C6018  ( .a(\prgm_register/n1957 ), .b(
        \prgm_register/n1958 ), .out(\prgm_register/or_signal [978]) );
  nand2 \prgm_register/C6019  ( .a(enable), .b(a[978]), .out(
        \prgm_register/n1959 ) );
  nand2 \prgm_register/C6020  ( .a(\prgm_register/en_not ), .b(a[979]), .out(
        \prgm_register/n1960 ) );
  nand2 \prgm_register/C6021  ( .a(\prgm_register/n1959 ), .b(
        \prgm_register/n1960 ), .out(\prgm_register/or_signal [979]) );
  nand2 \prgm_register/C6022  ( .a(enable), .b(a[979]), .out(
        \prgm_register/n1961 ) );
  nand2 \prgm_register/C6023  ( .a(\prgm_register/en_not ), .b(a[980]), .out(
        \prgm_register/n1962 ) );
  nand2 \prgm_register/C6024  ( .a(\prgm_register/n1961 ), .b(
        \prgm_register/n1962 ), .out(\prgm_register/or_signal [980]) );
  nand2 \prgm_register/C6025  ( .a(enable), .b(a[980]), .out(
        \prgm_register/n1963 ) );
  nand2 \prgm_register/C6026  ( .a(\prgm_register/en_not ), .b(a[981]), .out(
        \prgm_register/n1964 ) );
  nand2 \prgm_register/C6027  ( .a(\prgm_register/n1963 ), .b(
        \prgm_register/n1964 ), .out(\prgm_register/or_signal [981]) );
  nand2 \prgm_register/C6028  ( .a(enable), .b(a[981]), .out(
        \prgm_register/n1965 ) );
  nand2 \prgm_register/C6029  ( .a(\prgm_register/en_not ), .b(a[982]), .out(
        \prgm_register/n1966 ) );
  nand2 \prgm_register/C6030  ( .a(\prgm_register/n1965 ), .b(
        \prgm_register/n1966 ), .out(\prgm_register/or_signal [982]) );
  nand2 \prgm_register/C6031  ( .a(enable), .b(a[982]), .out(
        \prgm_register/n1967 ) );
  nand2 \prgm_register/C6032  ( .a(\prgm_register/en_not ), .b(a[983]), .out(
        \prgm_register/n1968 ) );
  nand2 \prgm_register/C6033  ( .a(\prgm_register/n1967 ), .b(
        \prgm_register/n1968 ), .out(\prgm_register/or_signal [983]) );
  nand2 \prgm_register/C6034  ( .a(enable), .b(a[983]), .out(
        \prgm_register/n1969 ) );
  nand2 \prgm_register/C6035  ( .a(\prgm_register/en_not ), .b(a[984]), .out(
        \prgm_register/n1970 ) );
  nand2 \prgm_register/C6036  ( .a(\prgm_register/n1969 ), .b(
        \prgm_register/n1970 ), .out(\prgm_register/or_signal [984]) );
  nand2 \prgm_register/C6037  ( .a(enable), .b(a[984]), .out(
        \prgm_register/n1971 ) );
  nand2 \prgm_register/C6038  ( .a(\prgm_register/en_not ), .b(a[985]), .out(
        \prgm_register/n1972 ) );
  nand2 \prgm_register/C6039  ( .a(\prgm_register/n1971 ), .b(
        \prgm_register/n1972 ), .out(\prgm_register/or_signal [985]) );
  nand2 \prgm_register/C6040  ( .a(enable), .b(a[985]), .out(
        \prgm_register/n1973 ) );
  nand2 \prgm_register/C6041  ( .a(\prgm_register/en_not ), .b(a[986]), .out(
        \prgm_register/n1974 ) );
  nand2 \prgm_register/C6042  ( .a(\prgm_register/n1973 ), .b(
        \prgm_register/n1974 ), .out(\prgm_register/or_signal [986]) );
  nand2 \prgm_register/C6043  ( .a(enable), .b(a[986]), .out(
        \prgm_register/n1975 ) );
  nand2 \prgm_register/C6044  ( .a(\prgm_register/en_not ), .b(a[987]), .out(
        \prgm_register/n1976 ) );
  nand2 \prgm_register/C6045  ( .a(\prgm_register/n1975 ), .b(
        \prgm_register/n1976 ), .out(\prgm_register/or_signal [987]) );
  nand2 \prgm_register/C6046  ( .a(enable), .b(a[987]), .out(
        \prgm_register/n1977 ) );
  nand2 \prgm_register/C6047  ( .a(\prgm_register/en_not ), .b(a[988]), .out(
        \prgm_register/n1978 ) );
  nand2 \prgm_register/C6048  ( .a(\prgm_register/n1977 ), .b(
        \prgm_register/n1978 ), .out(\prgm_register/or_signal [988]) );
  nand2 \prgm_register/C6049  ( .a(enable), .b(a[988]), .out(
        \prgm_register/n1979 ) );
  nand2 \prgm_register/C6050  ( .a(\prgm_register/en_not ), .b(a[989]), .out(
        \prgm_register/n1980 ) );
  nand2 \prgm_register/C6051  ( .a(\prgm_register/n1979 ), .b(
        \prgm_register/n1980 ), .out(\prgm_register/or_signal [989]) );
  nand2 \prgm_register/C6052  ( .a(enable), .b(a[989]), .out(
        \prgm_register/n1981 ) );
  nand2 \prgm_register/C6053  ( .a(\prgm_register/en_not ), .b(a[990]), .out(
        \prgm_register/n1982 ) );
  nand2 \prgm_register/C6054  ( .a(\prgm_register/n1981 ), .b(
        \prgm_register/n1982 ), .out(\prgm_register/or_signal [990]) );
  nand2 \prgm_register/C6055  ( .a(enable), .b(a[990]), .out(
        \prgm_register/n1983 ) );
  nand2 \prgm_register/C6056  ( .a(\prgm_register/en_not ), .b(a[991]), .out(
        \prgm_register/n1984 ) );
  nand2 \prgm_register/C6057  ( .a(\prgm_register/n1983 ), .b(
        \prgm_register/n1984 ), .out(\prgm_register/or_signal [991]) );
  nand2 \prgm_register/C6058  ( .a(enable), .b(a[991]), .out(
        \prgm_register/n1985 ) );
  nand2 \prgm_register/C6059  ( .a(\prgm_register/en_not ), .b(a[992]), .out(
        \prgm_register/n1986 ) );
  nand2 \prgm_register/C6060  ( .a(\prgm_register/n1985 ), .b(
        \prgm_register/n1986 ), .out(\prgm_register/or_signal [992]) );
  nand2 \prgm_register/C6061  ( .a(enable), .b(a[992]), .out(
        \prgm_register/n1987 ) );
  nand2 \prgm_register/C6062  ( .a(\prgm_register/en_not ), .b(a[993]), .out(
        \prgm_register/n1988 ) );
  nand2 \prgm_register/C6063  ( .a(\prgm_register/n1987 ), .b(
        \prgm_register/n1988 ), .out(\prgm_register/or_signal [993]) );
  nand2 \prgm_register/C6064  ( .a(enable), .b(a[993]), .out(
        \prgm_register/n1989 ) );
  nand2 \prgm_register/C6065  ( .a(\prgm_register/en_not ), .b(a[994]), .out(
        \prgm_register/n1990 ) );
  nand2 \prgm_register/C6066  ( .a(\prgm_register/n1989 ), .b(
        \prgm_register/n1990 ), .out(\prgm_register/or_signal [994]) );
  nand2 \prgm_register/C6067  ( .a(enable), .b(a[994]), .out(
        \prgm_register/n1991 ) );
  nand2 \prgm_register/C6068  ( .a(\prgm_register/en_not ), .b(a[995]), .out(
        \prgm_register/n1992 ) );
  nand2 \prgm_register/C6069  ( .a(\prgm_register/n1991 ), .b(
        \prgm_register/n1992 ), .out(\prgm_register/or_signal [995]) );
  nand2 \prgm_register/C6070  ( .a(enable), .b(a[995]), .out(
        \prgm_register/n1993 ) );
  nand2 \prgm_register/C6071  ( .a(\prgm_register/en_not ), .b(a[996]), .out(
        \prgm_register/n1994 ) );
  nand2 \prgm_register/C6072  ( .a(\prgm_register/n1993 ), .b(
        \prgm_register/n1994 ), .out(\prgm_register/or_signal [996]) );
  nand2 \prgm_register/C6073  ( .a(enable), .b(a[996]), .out(
        \prgm_register/n1995 ) );
  nand2 \prgm_register/C6074  ( .a(\prgm_register/en_not ), .b(a[997]), .out(
        \prgm_register/n1996 ) );
  nand2 \prgm_register/C6075  ( .a(\prgm_register/n1995 ), .b(
        \prgm_register/n1996 ), .out(\prgm_register/or_signal [997]) );
  nand2 \prgm_register/C6076  ( .a(enable), .b(a[997]), .out(
        \prgm_register/n1997 ) );
  nand2 \prgm_register/C6077  ( .a(\prgm_register/en_not ), .b(a[998]), .out(
        \prgm_register/n1998 ) );
  nand2 \prgm_register/C6078  ( .a(\prgm_register/n1997 ), .b(
        \prgm_register/n1998 ), .out(\prgm_register/or_signal [998]) );
  nand2 \prgm_register/C6079  ( .a(enable), .b(a[998]), .out(
        \prgm_register/n1999 ) );
  nand2 \prgm_register/C6080  ( .a(\prgm_register/en_not ), .b(a[999]), .out(
        \prgm_register/n2000 ) );
  nand2 \prgm_register/C6081  ( .a(\prgm_register/n1999 ), .b(
        \prgm_register/n2000 ), .out(\prgm_register/or_signal [999]) );
  nand2 \prgm_register/C6082  ( .a(enable), .b(a[999]), .out(
        \prgm_register/n2001 ) );
  nand2 \prgm_register/C6083  ( .a(\prgm_register/en_not ), .b(a[1000]), .out(
        \prgm_register/n2002 ) );
  nand2 \prgm_register/C6084  ( .a(\prgm_register/n2001 ), .b(
        \prgm_register/n2002 ), .out(\prgm_register/or_signal [1000]) );
  nand2 \prgm_register/C6085  ( .a(enable), .b(a[1000]), .out(
        \prgm_register/n2003 ) );
  nand2 \prgm_register/C6086  ( .a(\prgm_register/en_not ), .b(a[1001]), .out(
        \prgm_register/n2004 ) );
  nand2 \prgm_register/C6087  ( .a(\prgm_register/n2003 ), .b(
        \prgm_register/n2004 ), .out(\prgm_register/or_signal [1001]) );
  nand2 \prgm_register/C6088  ( .a(enable), .b(a[1001]), .out(
        \prgm_register/n2005 ) );
  nand2 \prgm_register/C6089  ( .a(\prgm_register/en_not ), .b(a[1002]), .out(
        \prgm_register/n2006 ) );
  nand2 \prgm_register/C6090  ( .a(\prgm_register/n2005 ), .b(
        \prgm_register/n2006 ), .out(\prgm_register/or_signal [1002]) );
  nand2 \prgm_register/C6091  ( .a(enable), .b(a[1002]), .out(
        \prgm_register/n2007 ) );
  nand2 \prgm_register/C6092  ( .a(\prgm_register/en_not ), .b(a[1003]), .out(
        \prgm_register/n2008 ) );
  nand2 \prgm_register/C6093  ( .a(\prgm_register/n2007 ), .b(
        \prgm_register/n2008 ), .out(\prgm_register/or_signal [1003]) );
  nand2 \prgm_register/C6094  ( .a(enable), .b(a[1003]), .out(
        \prgm_register/n2009 ) );
  nand2 \prgm_register/C6095  ( .a(\prgm_register/en_not ), .b(a[1004]), .out(
        \prgm_register/n2010 ) );
  nand2 \prgm_register/C6096  ( .a(\prgm_register/n2009 ), .b(
        \prgm_register/n2010 ), .out(\prgm_register/or_signal [1004]) );
  nand2 \prgm_register/C6097  ( .a(enable), .b(a[1004]), .out(
        \prgm_register/n2011 ) );
  nand2 \prgm_register/C6098  ( .a(\prgm_register/en_not ), .b(a[1005]), .out(
        \prgm_register/n2012 ) );
  nand2 \prgm_register/C6099  ( .a(\prgm_register/n2011 ), .b(
        \prgm_register/n2012 ), .out(\prgm_register/or_signal [1005]) );
  nand2 \prgm_register/C6100  ( .a(enable), .b(a[1005]), .out(
        \prgm_register/n2013 ) );
  nand2 \prgm_register/C6101  ( .a(\prgm_register/en_not ), .b(a[1006]), .out(
        \prgm_register/n2014 ) );
  nand2 \prgm_register/C6102  ( .a(\prgm_register/n2013 ), .b(
        \prgm_register/n2014 ), .out(\prgm_register/or_signal [1006]) );
  nand2 \prgm_register/C6103  ( .a(enable), .b(a[1006]), .out(
        \prgm_register/n2015 ) );
  nand2 \prgm_register/C6104  ( .a(\prgm_register/en_not ), .b(a[1007]), .out(
        \prgm_register/n2016 ) );
  nand2 \prgm_register/C6105  ( .a(\prgm_register/n2015 ), .b(
        \prgm_register/n2016 ), .out(\prgm_register/or_signal [1007]) );
  nand2 \prgm_register/C6106  ( .a(enable), .b(a[1007]), .out(
        \prgm_register/n2017 ) );
  nand2 \prgm_register/C6107  ( .a(\prgm_register/en_not ), .b(a[1008]), .out(
        \prgm_register/n2018 ) );
  nand2 \prgm_register/C6108  ( .a(\prgm_register/n2017 ), .b(
        \prgm_register/n2018 ), .out(\prgm_register/or_signal [1008]) );
  nand2 \prgm_register/C6109  ( .a(enable), .b(a[1008]), .out(
        \prgm_register/n2019 ) );
  nand2 \prgm_register/C6110  ( .a(\prgm_register/en_not ), .b(a[1009]), .out(
        \prgm_register/n2020 ) );
  nand2 \prgm_register/C6111  ( .a(\prgm_register/n2019 ), .b(
        \prgm_register/n2020 ), .out(\prgm_register/or_signal [1009]) );
  nand2 \prgm_register/C6112  ( .a(enable), .b(a[1009]), .out(
        \prgm_register/n2021 ) );
  nand2 \prgm_register/C6113  ( .a(\prgm_register/en_not ), .b(a[1010]), .out(
        \prgm_register/n2022 ) );
  nand2 \prgm_register/C6114  ( .a(\prgm_register/n2021 ), .b(
        \prgm_register/n2022 ), .out(\prgm_register/or_signal [1010]) );
  nand2 \prgm_register/C6115  ( .a(enable), .b(a[1010]), .out(
        \prgm_register/n2023 ) );
  nand2 \prgm_register/C6116  ( .a(\prgm_register/en_not ), .b(a[1011]), .out(
        \prgm_register/n2024 ) );
  nand2 \prgm_register/C6117  ( .a(\prgm_register/n2023 ), .b(
        \prgm_register/n2024 ), .out(\prgm_register/or_signal [1011]) );
  nand2 \prgm_register/C6118  ( .a(enable), .b(a[1011]), .out(
        \prgm_register/n2025 ) );
  nand2 \prgm_register/C6119  ( .a(\prgm_register/en_not ), .b(a[1012]), .out(
        \prgm_register/n2026 ) );
  nand2 \prgm_register/C6120  ( .a(\prgm_register/n2025 ), .b(
        \prgm_register/n2026 ), .out(\prgm_register/or_signal [1012]) );
  nand2 \prgm_register/C6121  ( .a(enable), .b(a[1012]), .out(
        \prgm_register/n2027 ) );
  nand2 \prgm_register/C6122  ( .a(\prgm_register/en_not ), .b(a[1013]), .out(
        \prgm_register/n2028 ) );
  nand2 \prgm_register/C6123  ( .a(\prgm_register/n2027 ), .b(
        \prgm_register/n2028 ), .out(\prgm_register/or_signal [1013]) );
  nand2 \prgm_register/C6124  ( .a(enable), .b(a[1013]), .out(
        \prgm_register/n2029 ) );
  nand2 \prgm_register/C6125  ( .a(\prgm_register/en_not ), .b(a[1014]), .out(
        \prgm_register/n2030 ) );
  nand2 \prgm_register/C6126  ( .a(\prgm_register/n2029 ), .b(
        \prgm_register/n2030 ), .out(\prgm_register/or_signal [1014]) );
  nand2 \prgm_register/C6127  ( .a(enable), .b(a[1014]), .out(
        \prgm_register/n2031 ) );
  nand2 \prgm_register/C6128  ( .a(\prgm_register/en_not ), .b(a[1015]), .out(
        \prgm_register/n2032 ) );
  nand2 \prgm_register/C6129  ( .a(\prgm_register/n2031 ), .b(
        \prgm_register/n2032 ), .out(\prgm_register/or_signal [1015]) );
  nand2 \prgm_register/C6130  ( .a(enable), .b(a[1015]), .out(
        \prgm_register/n2033 ) );
  nand2 \prgm_register/C6131  ( .a(\prgm_register/en_not ), .b(a[1016]), .out(
        \prgm_register/n2034 ) );
  nand2 \prgm_register/C6132  ( .a(\prgm_register/n2033 ), .b(
        \prgm_register/n2034 ), .out(\prgm_register/or_signal [1016]) );
  nand2 \prgm_register/C6133  ( .a(enable), .b(a[1016]), .out(
        \prgm_register/n2035 ) );
  nand2 \prgm_register/C6134  ( .a(\prgm_register/en_not ), .b(a[1017]), .out(
        \prgm_register/n2036 ) );
  nand2 \prgm_register/C6135  ( .a(\prgm_register/n2035 ), .b(
        \prgm_register/n2036 ), .out(\prgm_register/or_signal [1017]) );
  nand2 \prgm_register/C6136  ( .a(enable), .b(a[1017]), .out(
        \prgm_register/n2037 ) );
  nand2 \prgm_register/C6137  ( .a(\prgm_register/en_not ), .b(a[1018]), .out(
        \prgm_register/n2038 ) );
  nand2 \prgm_register/C6138  ( .a(\prgm_register/n2037 ), .b(
        \prgm_register/n2038 ), .out(\prgm_register/or_signal [1018]) );
  nand2 \prgm_register/C6139  ( .a(enable), .b(a[1018]), .out(
        \prgm_register/n2039 ) );
  nand2 \prgm_register/C6140  ( .a(\prgm_register/en_not ), .b(a[1019]), .out(
        \prgm_register/n2040 ) );
  nand2 \prgm_register/C6141  ( .a(\prgm_register/n2039 ), .b(
        \prgm_register/n2040 ), .out(\prgm_register/or_signal [1019]) );
  nand2 \prgm_register/C6142  ( .a(enable), .b(a[1019]), .out(
        \prgm_register/n2041 ) );
  nand2 \prgm_register/C6143  ( .a(\prgm_register/en_not ), .b(a[1020]), .out(
        \prgm_register/n2042 ) );
  nand2 \prgm_register/C6144  ( .a(\prgm_register/n2041 ), .b(
        \prgm_register/n2042 ), .out(\prgm_register/or_signal [1020]) );
  nand2 \prgm_register/C6145  ( .a(enable), .b(a[1020]), .out(
        \prgm_register/n2043 ) );
  nand2 \prgm_register/C6146  ( .a(\prgm_register/en_not ), .b(a[1021]), .out(
        \prgm_register/n2044 ) );
  nand2 \prgm_register/C6147  ( .a(\prgm_register/n2043 ), .b(
        \prgm_register/n2044 ), .out(\prgm_register/or_signal [1021]) );
  nand2 \prgm_register/C6148  ( .a(enable), .b(a[1021]), .out(
        \prgm_register/n2045 ) );
  nand2 \prgm_register/C6149  ( .a(\prgm_register/en_not ), .b(a[1022]), .out(
        \prgm_register/n2046 ) );
  nand2 \prgm_register/C6150  ( .a(\prgm_register/n2045 ), .b(
        \prgm_register/n2046 ), .out(\prgm_register/or_signal [1022]) );
  nand2 \prgm_register/C6151  ( .a(enable), .b(a[1022]), .out(
        \prgm_register/n2047 ) );
  nand2 \prgm_register/C6152  ( .a(\prgm_register/en_not ), .b(a[1023]), .out(
        \prgm_register/n2048 ) );
  nand2 \prgm_register/C6153  ( .a(\prgm_register/n2047 ), .b(
        \prgm_register/n2048 ), .out(\prgm_register/or_signal [1023]) );
  d_ff \prgm_register/genblk1[1023].single_DFF  ( .d(
        \prgm_register/or_signal [1023]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1023]) );
  d_ff \prgm_register/genblk1[1022].single_DFF  ( .d(
        \prgm_register/or_signal [1022]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1022]) );
  d_ff \prgm_register/genblk1[1021].single_DFF  ( .d(
        \prgm_register/or_signal [1021]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1021]) );
  d_ff \prgm_register/genblk1[1020].single_DFF  ( .d(
        \prgm_register/or_signal [1020]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1020]) );
  d_ff \prgm_register/genblk1[1019].single_DFF  ( .d(
        \prgm_register/or_signal [1019]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1019]) );
  d_ff \prgm_register/genblk1[1018].single_DFF  ( .d(
        \prgm_register/or_signal [1018]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1018]) );
  d_ff \prgm_register/genblk1[1017].single_DFF  ( .d(
        \prgm_register/or_signal [1017]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1017]) );
  d_ff \prgm_register/genblk1[1016].single_DFF  ( .d(
        \prgm_register/or_signal [1016]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1016]) );
  d_ff \prgm_register/genblk1[1015].single_DFF  ( .d(
        \prgm_register/or_signal [1015]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1015]) );
  d_ff \prgm_register/genblk1[1014].single_DFF  ( .d(
        \prgm_register/or_signal [1014]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1014]) );
  d_ff \prgm_register/genblk1[1013].single_DFF  ( .d(
        \prgm_register/or_signal [1013]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1013]) );
  d_ff \prgm_register/genblk1[1012].single_DFF  ( .d(
        \prgm_register/or_signal [1012]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1012]) );
  d_ff \prgm_register/genblk1[1011].single_DFF  ( .d(
        \prgm_register/or_signal [1011]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1011]) );
  d_ff \prgm_register/genblk1[1010].single_DFF  ( .d(
        \prgm_register/or_signal [1010]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1010]) );
  d_ff \prgm_register/genblk1[1009].single_DFF  ( .d(
        \prgm_register/or_signal [1009]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1009]) );
  d_ff \prgm_register/genblk1[1008].single_DFF  ( .d(
        \prgm_register/or_signal [1008]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1008]) );
  d_ff \prgm_register/genblk1[1007].single_DFF  ( .d(
        \prgm_register/or_signal [1007]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1007]) );
  d_ff \prgm_register/genblk1[1006].single_DFF  ( .d(
        \prgm_register/or_signal [1006]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1006]) );
  d_ff \prgm_register/genblk1[1005].single_DFF  ( .d(
        \prgm_register/or_signal [1005]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1005]) );
  d_ff \prgm_register/genblk1[1004].single_DFF  ( .d(
        \prgm_register/or_signal [1004]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1004]) );
  d_ff \prgm_register/genblk1[1003].single_DFF  ( .d(
        \prgm_register/or_signal [1003]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1003]) );
  d_ff \prgm_register/genblk1[1002].single_DFF  ( .d(
        \prgm_register/or_signal [1002]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1002]) );
  d_ff \prgm_register/genblk1[1001].single_DFF  ( .d(
        \prgm_register/or_signal [1001]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1001]) );
  d_ff \prgm_register/genblk1[1000].single_DFF  ( .d(
        \prgm_register/or_signal [1000]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[1000]) );
  d_ff \prgm_register/genblk1[999].single_DFF  ( .d(
        \prgm_register/or_signal [999]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[999]) );
  d_ff \prgm_register/genblk1[998].single_DFF  ( .d(
        \prgm_register/or_signal [998]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[998]) );
  d_ff \prgm_register/genblk1[997].single_DFF  ( .d(
        \prgm_register/or_signal [997]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[997]) );
  d_ff \prgm_register/genblk1[996].single_DFF  ( .d(
        \prgm_register/or_signal [996]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[996]) );
  d_ff \prgm_register/genblk1[995].single_DFF  ( .d(
        \prgm_register/or_signal [995]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[995]) );
  d_ff \prgm_register/genblk1[994].single_DFF  ( .d(
        \prgm_register/or_signal [994]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[994]) );
  d_ff \prgm_register/genblk1[993].single_DFF  ( .d(
        \prgm_register/or_signal [993]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[993]) );
  d_ff \prgm_register/genblk1[992].single_DFF  ( .d(
        \prgm_register/or_signal [992]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[992]) );
  d_ff \prgm_register/genblk1[991].single_DFF  ( .d(
        \prgm_register/or_signal [991]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[991]) );
  d_ff \prgm_register/genblk1[990].single_DFF  ( .d(
        \prgm_register/or_signal [990]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[990]) );
  d_ff \prgm_register/genblk1[989].single_DFF  ( .d(
        \prgm_register/or_signal [989]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[989]) );
  d_ff \prgm_register/genblk1[988].single_DFF  ( .d(
        \prgm_register/or_signal [988]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[988]) );
  d_ff \prgm_register/genblk1[987].single_DFF  ( .d(
        \prgm_register/or_signal [987]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[987]) );
  d_ff \prgm_register/genblk1[986].single_DFF  ( .d(
        \prgm_register/or_signal [986]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[986]) );
  d_ff \prgm_register/genblk1[985].single_DFF  ( .d(
        \prgm_register/or_signal [985]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[985]) );
  d_ff \prgm_register/genblk1[984].single_DFF  ( .d(
        \prgm_register/or_signal [984]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[984]) );
  d_ff \prgm_register/genblk1[983].single_DFF  ( .d(
        \prgm_register/or_signal [983]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[983]) );
  d_ff \prgm_register/genblk1[982].single_DFF  ( .d(
        \prgm_register/or_signal [982]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[982]) );
  d_ff \prgm_register/genblk1[981].single_DFF  ( .d(
        \prgm_register/or_signal [981]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[981]) );
  d_ff \prgm_register/genblk1[980].single_DFF  ( .d(
        \prgm_register/or_signal [980]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[980]) );
  d_ff \prgm_register/genblk1[979].single_DFF  ( .d(
        \prgm_register/or_signal [979]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[979]) );
  d_ff \prgm_register/genblk1[978].single_DFF  ( .d(
        \prgm_register/or_signal [978]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[978]) );
  d_ff \prgm_register/genblk1[977].single_DFF  ( .d(
        \prgm_register/or_signal [977]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[977]) );
  d_ff \prgm_register/genblk1[976].single_DFF  ( .d(
        \prgm_register/or_signal [976]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[976]) );
  d_ff \prgm_register/genblk1[975].single_DFF  ( .d(
        \prgm_register/or_signal [975]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[975]) );
  d_ff \prgm_register/genblk1[974].single_DFF  ( .d(
        \prgm_register/or_signal [974]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[974]) );
  d_ff \prgm_register/genblk1[973].single_DFF  ( .d(
        \prgm_register/or_signal [973]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[973]) );
  d_ff \prgm_register/genblk1[972].single_DFF  ( .d(
        \prgm_register/or_signal [972]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[972]) );
  d_ff \prgm_register/genblk1[971].single_DFF  ( .d(
        \prgm_register/or_signal [971]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[971]) );
  d_ff \prgm_register/genblk1[970].single_DFF  ( .d(
        \prgm_register/or_signal [970]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[970]) );
  d_ff \prgm_register/genblk1[969].single_DFF  ( .d(
        \prgm_register/or_signal [969]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[969]) );
  d_ff \prgm_register/genblk1[968].single_DFF  ( .d(
        \prgm_register/or_signal [968]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[968]) );
  d_ff \prgm_register/genblk1[967].single_DFF  ( .d(
        \prgm_register/or_signal [967]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[967]) );
  d_ff \prgm_register/genblk1[966].single_DFF  ( .d(
        \prgm_register/or_signal [966]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[966]) );
  d_ff \prgm_register/genblk1[965].single_DFF  ( .d(
        \prgm_register/or_signal [965]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[965]) );
  d_ff \prgm_register/genblk1[964].single_DFF  ( .d(
        \prgm_register/or_signal [964]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[964]) );
  d_ff \prgm_register/genblk1[963].single_DFF  ( .d(
        \prgm_register/or_signal [963]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[963]) );
  d_ff \prgm_register/genblk1[962].single_DFF  ( .d(
        \prgm_register/or_signal [962]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[962]) );
  d_ff \prgm_register/genblk1[961].single_DFF  ( .d(
        \prgm_register/or_signal [961]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[961]) );
  d_ff \prgm_register/genblk1[960].single_DFF  ( .d(
        \prgm_register/or_signal [960]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[960]) );
  d_ff \prgm_register/genblk1[959].single_DFF  ( .d(
        \prgm_register/or_signal [959]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[959]) );
  d_ff \prgm_register/genblk1[958].single_DFF  ( .d(
        \prgm_register/or_signal [958]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[958]) );
  d_ff \prgm_register/genblk1[957].single_DFF  ( .d(
        \prgm_register/or_signal [957]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[957]) );
  d_ff \prgm_register/genblk1[956].single_DFF  ( .d(
        \prgm_register/or_signal [956]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[956]) );
  d_ff \prgm_register/genblk1[955].single_DFF  ( .d(
        \prgm_register/or_signal [955]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[955]) );
  d_ff \prgm_register/genblk1[954].single_DFF  ( .d(
        \prgm_register/or_signal [954]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[954]) );
  d_ff \prgm_register/genblk1[953].single_DFF  ( .d(
        \prgm_register/or_signal [953]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[953]) );
  d_ff \prgm_register/genblk1[952].single_DFF  ( .d(
        \prgm_register/or_signal [952]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[952]) );
  d_ff \prgm_register/genblk1[951].single_DFF  ( .d(
        \prgm_register/or_signal [951]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[951]) );
  d_ff \prgm_register/genblk1[950].single_DFF  ( .d(
        \prgm_register/or_signal [950]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[950]) );
  d_ff \prgm_register/genblk1[949].single_DFF  ( .d(
        \prgm_register/or_signal [949]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[949]) );
  d_ff \prgm_register/genblk1[948].single_DFF  ( .d(
        \prgm_register/or_signal [948]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[948]) );
  d_ff \prgm_register/genblk1[947].single_DFF  ( .d(
        \prgm_register/or_signal [947]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[947]) );
  d_ff \prgm_register/genblk1[946].single_DFF  ( .d(
        \prgm_register/or_signal [946]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[946]) );
  d_ff \prgm_register/genblk1[945].single_DFF  ( .d(
        \prgm_register/or_signal [945]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[945]) );
  d_ff \prgm_register/genblk1[944].single_DFF  ( .d(
        \prgm_register/or_signal [944]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[944]) );
  d_ff \prgm_register/genblk1[943].single_DFF  ( .d(
        \prgm_register/or_signal [943]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[943]) );
  d_ff \prgm_register/genblk1[942].single_DFF  ( .d(
        \prgm_register/or_signal [942]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[942]) );
  d_ff \prgm_register/genblk1[941].single_DFF  ( .d(
        \prgm_register/or_signal [941]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[941]) );
  d_ff \prgm_register/genblk1[940].single_DFF  ( .d(
        \prgm_register/or_signal [940]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[940]) );
  d_ff \prgm_register/genblk1[939].single_DFF  ( .d(
        \prgm_register/or_signal [939]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[939]) );
  d_ff \prgm_register/genblk1[938].single_DFF  ( .d(
        \prgm_register/or_signal [938]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[938]) );
  d_ff \prgm_register/genblk1[937].single_DFF  ( .d(
        \prgm_register/or_signal [937]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[937]) );
  d_ff \prgm_register/genblk1[936].single_DFF  ( .d(
        \prgm_register/or_signal [936]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[936]) );
  d_ff \prgm_register/genblk1[935].single_DFF  ( .d(
        \prgm_register/or_signal [935]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[935]) );
  d_ff \prgm_register/genblk1[934].single_DFF  ( .d(
        \prgm_register/or_signal [934]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[934]) );
  d_ff \prgm_register/genblk1[933].single_DFF  ( .d(
        \prgm_register/or_signal [933]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[933]) );
  d_ff \prgm_register/genblk1[932].single_DFF  ( .d(
        \prgm_register/or_signal [932]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[932]) );
  d_ff \prgm_register/genblk1[931].single_DFF  ( .d(
        \prgm_register/or_signal [931]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[931]) );
  d_ff \prgm_register/genblk1[930].single_DFF  ( .d(
        \prgm_register/or_signal [930]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[930]) );
  d_ff \prgm_register/genblk1[929].single_DFF  ( .d(
        \prgm_register/or_signal [929]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[929]) );
  d_ff \prgm_register/genblk1[928].single_DFF  ( .d(
        \prgm_register/or_signal [928]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[928]) );
  d_ff \prgm_register/genblk1[927].single_DFF  ( .d(
        \prgm_register/or_signal [927]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[927]) );
  d_ff \prgm_register/genblk1[926].single_DFF  ( .d(
        \prgm_register/or_signal [926]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[926]) );
  d_ff \prgm_register/genblk1[925].single_DFF  ( .d(
        \prgm_register/or_signal [925]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[925]) );
  d_ff \prgm_register/genblk1[924].single_DFF  ( .d(
        \prgm_register/or_signal [924]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[924]) );
  d_ff \prgm_register/genblk1[923].single_DFF  ( .d(
        \prgm_register/or_signal [923]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[923]) );
  d_ff \prgm_register/genblk1[922].single_DFF  ( .d(
        \prgm_register/or_signal [922]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[922]) );
  d_ff \prgm_register/genblk1[921].single_DFF  ( .d(
        \prgm_register/or_signal [921]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[921]) );
  d_ff \prgm_register/genblk1[920].single_DFF  ( .d(
        \prgm_register/or_signal [920]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[920]) );
  d_ff \prgm_register/genblk1[919].single_DFF  ( .d(
        \prgm_register/or_signal [919]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[919]) );
  d_ff \prgm_register/genblk1[918].single_DFF  ( .d(
        \prgm_register/or_signal [918]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[918]) );
  d_ff \prgm_register/genblk1[917].single_DFF  ( .d(
        \prgm_register/or_signal [917]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[917]) );
  d_ff \prgm_register/genblk1[916].single_DFF  ( .d(
        \prgm_register/or_signal [916]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[916]) );
  d_ff \prgm_register/genblk1[915].single_DFF  ( .d(
        \prgm_register/or_signal [915]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[915]) );
  d_ff \prgm_register/genblk1[914].single_DFF  ( .d(
        \prgm_register/or_signal [914]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[914]) );
  d_ff \prgm_register/genblk1[913].single_DFF  ( .d(
        \prgm_register/or_signal [913]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[913]) );
  d_ff \prgm_register/genblk1[912].single_DFF  ( .d(
        \prgm_register/or_signal [912]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[912]) );
  d_ff \prgm_register/genblk1[911].single_DFF  ( .d(
        \prgm_register/or_signal [911]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[911]) );
  d_ff \prgm_register/genblk1[910].single_DFF  ( .d(
        \prgm_register/or_signal [910]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[910]) );
  d_ff \prgm_register/genblk1[909].single_DFF  ( .d(
        \prgm_register/or_signal [909]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[909]) );
  d_ff \prgm_register/genblk1[908].single_DFF  ( .d(
        \prgm_register/or_signal [908]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[908]) );
  d_ff \prgm_register/genblk1[907].single_DFF  ( .d(
        \prgm_register/or_signal [907]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[907]) );
  d_ff \prgm_register/genblk1[906].single_DFF  ( .d(
        \prgm_register/or_signal [906]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[906]) );
  d_ff \prgm_register/genblk1[905].single_DFF  ( .d(
        \prgm_register/or_signal [905]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[905]) );
  d_ff \prgm_register/genblk1[904].single_DFF  ( .d(
        \prgm_register/or_signal [904]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[904]) );
  d_ff \prgm_register/genblk1[903].single_DFF  ( .d(
        \prgm_register/or_signal [903]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[903]) );
  d_ff \prgm_register/genblk1[902].single_DFF  ( .d(
        \prgm_register/or_signal [902]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[902]) );
  d_ff \prgm_register/genblk1[901].single_DFF  ( .d(
        \prgm_register/or_signal [901]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[901]) );
  d_ff \prgm_register/genblk1[900].single_DFF  ( .d(
        \prgm_register/or_signal [900]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[900]) );
  d_ff \prgm_register/genblk1[899].single_DFF  ( .d(
        \prgm_register/or_signal [899]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[899]) );
  d_ff \prgm_register/genblk1[898].single_DFF  ( .d(
        \prgm_register/or_signal [898]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[898]) );
  d_ff \prgm_register/genblk1[897].single_DFF  ( .d(
        \prgm_register/or_signal [897]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[897]) );
  d_ff \prgm_register/genblk1[896].single_DFF  ( .d(
        \prgm_register/or_signal [896]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[896]) );
  d_ff \prgm_register/genblk1[895].single_DFF  ( .d(
        \prgm_register/or_signal [895]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[895]) );
  d_ff \prgm_register/genblk1[894].single_DFF  ( .d(
        \prgm_register/or_signal [894]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[894]) );
  d_ff \prgm_register/genblk1[893].single_DFF  ( .d(
        \prgm_register/or_signal [893]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[893]) );
  d_ff \prgm_register/genblk1[892].single_DFF  ( .d(
        \prgm_register/or_signal [892]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[892]) );
  d_ff \prgm_register/genblk1[891].single_DFF  ( .d(
        \prgm_register/or_signal [891]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[891]) );
  d_ff \prgm_register/genblk1[890].single_DFF  ( .d(
        \prgm_register/or_signal [890]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[890]) );
  d_ff \prgm_register/genblk1[889].single_DFF  ( .d(
        \prgm_register/or_signal [889]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[889]) );
  d_ff \prgm_register/genblk1[888].single_DFF  ( .d(
        \prgm_register/or_signal [888]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[888]) );
  d_ff \prgm_register/genblk1[887].single_DFF  ( .d(
        \prgm_register/or_signal [887]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[887]) );
  d_ff \prgm_register/genblk1[886].single_DFF  ( .d(
        \prgm_register/or_signal [886]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[886]) );
  d_ff \prgm_register/genblk1[885].single_DFF  ( .d(
        \prgm_register/or_signal [885]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[885]) );
  d_ff \prgm_register/genblk1[884].single_DFF  ( .d(
        \prgm_register/or_signal [884]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[884]) );
  d_ff \prgm_register/genblk1[883].single_DFF  ( .d(
        \prgm_register/or_signal [883]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[883]) );
  d_ff \prgm_register/genblk1[882].single_DFF  ( .d(
        \prgm_register/or_signal [882]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[882]) );
  d_ff \prgm_register/genblk1[881].single_DFF  ( .d(
        \prgm_register/or_signal [881]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[881]) );
  d_ff \prgm_register/genblk1[880].single_DFF  ( .d(
        \prgm_register/or_signal [880]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[880]) );
  d_ff \prgm_register/genblk1[879].single_DFF  ( .d(
        \prgm_register/or_signal [879]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[879]) );
  d_ff \prgm_register/genblk1[878].single_DFF  ( .d(
        \prgm_register/or_signal [878]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[878]) );
  d_ff \prgm_register/genblk1[877].single_DFF  ( .d(
        \prgm_register/or_signal [877]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[877]) );
  d_ff \prgm_register/genblk1[876].single_DFF  ( .d(
        \prgm_register/or_signal [876]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[876]) );
  d_ff \prgm_register/genblk1[875].single_DFF  ( .d(
        \prgm_register/or_signal [875]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[875]) );
  d_ff \prgm_register/genblk1[874].single_DFF  ( .d(
        \prgm_register/or_signal [874]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[874]) );
  d_ff \prgm_register/genblk1[873].single_DFF  ( .d(
        \prgm_register/or_signal [873]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[873]) );
  d_ff \prgm_register/genblk1[872].single_DFF  ( .d(
        \prgm_register/or_signal [872]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[872]) );
  d_ff \prgm_register/genblk1[871].single_DFF  ( .d(
        \prgm_register/or_signal [871]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[871]) );
  d_ff \prgm_register/genblk1[870].single_DFF  ( .d(
        \prgm_register/or_signal [870]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[870]) );
  d_ff \prgm_register/genblk1[869].single_DFF  ( .d(
        \prgm_register/or_signal [869]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[869]) );
  d_ff \prgm_register/genblk1[868].single_DFF  ( .d(
        \prgm_register/or_signal [868]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[868]) );
  d_ff \prgm_register/genblk1[867].single_DFF  ( .d(
        \prgm_register/or_signal [867]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[867]) );
  d_ff \prgm_register/genblk1[866].single_DFF  ( .d(
        \prgm_register/or_signal [866]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[866]) );
  d_ff \prgm_register/genblk1[865].single_DFF  ( .d(
        \prgm_register/or_signal [865]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[865]) );
  d_ff \prgm_register/genblk1[864].single_DFF  ( .d(
        \prgm_register/or_signal [864]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[864]) );
  d_ff \prgm_register/genblk1[863].single_DFF  ( .d(
        \prgm_register/or_signal [863]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[863]) );
  d_ff \prgm_register/genblk1[862].single_DFF  ( .d(
        \prgm_register/or_signal [862]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[862]) );
  d_ff \prgm_register/genblk1[861].single_DFF  ( .d(
        \prgm_register/or_signal [861]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[861]) );
  d_ff \prgm_register/genblk1[860].single_DFF  ( .d(
        \prgm_register/or_signal [860]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[860]) );
  d_ff \prgm_register/genblk1[859].single_DFF  ( .d(
        \prgm_register/or_signal [859]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[859]) );
  d_ff \prgm_register/genblk1[858].single_DFF  ( .d(
        \prgm_register/or_signal [858]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[858]) );
  d_ff \prgm_register/genblk1[857].single_DFF  ( .d(
        \prgm_register/or_signal [857]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[857]) );
  d_ff \prgm_register/genblk1[856].single_DFF  ( .d(
        \prgm_register/or_signal [856]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[856]) );
  d_ff \prgm_register/genblk1[855].single_DFF  ( .d(
        \prgm_register/or_signal [855]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[855]) );
  d_ff \prgm_register/genblk1[854].single_DFF  ( .d(
        \prgm_register/or_signal [854]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[854]) );
  d_ff \prgm_register/genblk1[853].single_DFF  ( .d(
        \prgm_register/or_signal [853]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[853]) );
  d_ff \prgm_register/genblk1[852].single_DFF  ( .d(
        \prgm_register/or_signal [852]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[852]) );
  d_ff \prgm_register/genblk1[851].single_DFF  ( .d(
        \prgm_register/or_signal [851]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[851]) );
  d_ff \prgm_register/genblk1[850].single_DFF  ( .d(
        \prgm_register/or_signal [850]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[850]) );
  d_ff \prgm_register/genblk1[849].single_DFF  ( .d(
        \prgm_register/or_signal [849]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[849]) );
  d_ff \prgm_register/genblk1[848].single_DFF  ( .d(
        \prgm_register/or_signal [848]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[848]) );
  d_ff \prgm_register/genblk1[847].single_DFF  ( .d(
        \prgm_register/or_signal [847]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[847]) );
  d_ff \prgm_register/genblk1[846].single_DFF  ( .d(
        \prgm_register/or_signal [846]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[846]) );
  d_ff \prgm_register/genblk1[845].single_DFF  ( .d(
        \prgm_register/or_signal [845]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[845]) );
  d_ff \prgm_register/genblk1[844].single_DFF  ( .d(
        \prgm_register/or_signal [844]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[844]) );
  d_ff \prgm_register/genblk1[843].single_DFF  ( .d(
        \prgm_register/or_signal [843]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[843]) );
  d_ff \prgm_register/genblk1[842].single_DFF  ( .d(
        \prgm_register/or_signal [842]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[842]) );
  d_ff \prgm_register/genblk1[841].single_DFF  ( .d(
        \prgm_register/or_signal [841]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[841]) );
  d_ff \prgm_register/genblk1[840].single_DFF  ( .d(
        \prgm_register/or_signal [840]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[840]) );
  d_ff \prgm_register/genblk1[839].single_DFF  ( .d(
        \prgm_register/or_signal [839]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[839]) );
  d_ff \prgm_register/genblk1[838].single_DFF  ( .d(
        \prgm_register/or_signal [838]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[838]) );
  d_ff \prgm_register/genblk1[837].single_DFF  ( .d(
        \prgm_register/or_signal [837]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[837]) );
  d_ff \prgm_register/genblk1[836].single_DFF  ( .d(
        \prgm_register/or_signal [836]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[836]) );
  d_ff \prgm_register/genblk1[835].single_DFF  ( .d(
        \prgm_register/or_signal [835]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[835]) );
  d_ff \prgm_register/genblk1[834].single_DFF  ( .d(
        \prgm_register/or_signal [834]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[834]) );
  d_ff \prgm_register/genblk1[833].single_DFF  ( .d(
        \prgm_register/or_signal [833]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[833]) );
  d_ff \prgm_register/genblk1[832].single_DFF  ( .d(
        \prgm_register/or_signal [832]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[832]) );
  d_ff \prgm_register/genblk1[831].single_DFF  ( .d(
        \prgm_register/or_signal [831]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[831]) );
  d_ff \prgm_register/genblk1[830].single_DFF  ( .d(
        \prgm_register/or_signal [830]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[830]) );
  d_ff \prgm_register/genblk1[829].single_DFF  ( .d(
        \prgm_register/or_signal [829]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[829]) );
  d_ff \prgm_register/genblk1[828].single_DFF  ( .d(
        \prgm_register/or_signal [828]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[828]) );
  d_ff \prgm_register/genblk1[827].single_DFF  ( .d(
        \prgm_register/or_signal [827]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[827]) );
  d_ff \prgm_register/genblk1[826].single_DFF  ( .d(
        \prgm_register/or_signal [826]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[826]) );
  d_ff \prgm_register/genblk1[825].single_DFF  ( .d(
        \prgm_register/or_signal [825]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[825]) );
  d_ff \prgm_register/genblk1[824].single_DFF  ( .d(
        \prgm_register/or_signal [824]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[824]) );
  d_ff \prgm_register/genblk1[823].single_DFF  ( .d(
        \prgm_register/or_signal [823]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[823]) );
  d_ff \prgm_register/genblk1[822].single_DFF  ( .d(
        \prgm_register/or_signal [822]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[822]) );
  d_ff \prgm_register/genblk1[821].single_DFF  ( .d(
        \prgm_register/or_signal [821]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[821]) );
  d_ff \prgm_register/genblk1[820].single_DFF  ( .d(
        \prgm_register/or_signal [820]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[820]) );
  d_ff \prgm_register/genblk1[819].single_DFF  ( .d(
        \prgm_register/or_signal [819]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[819]) );
  d_ff \prgm_register/genblk1[818].single_DFF  ( .d(
        \prgm_register/or_signal [818]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[818]) );
  d_ff \prgm_register/genblk1[817].single_DFF  ( .d(
        \prgm_register/or_signal [817]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[817]) );
  d_ff \prgm_register/genblk1[816].single_DFF  ( .d(
        \prgm_register/or_signal [816]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[816]) );
  d_ff \prgm_register/genblk1[815].single_DFF  ( .d(
        \prgm_register/or_signal [815]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[815]) );
  d_ff \prgm_register/genblk1[814].single_DFF  ( .d(
        \prgm_register/or_signal [814]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[814]) );
  d_ff \prgm_register/genblk1[813].single_DFF  ( .d(
        \prgm_register/or_signal [813]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[813]) );
  d_ff \prgm_register/genblk1[812].single_DFF  ( .d(
        \prgm_register/or_signal [812]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[812]) );
  d_ff \prgm_register/genblk1[811].single_DFF  ( .d(
        \prgm_register/or_signal [811]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[811]) );
  d_ff \prgm_register/genblk1[810].single_DFF  ( .d(
        \prgm_register/or_signal [810]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[810]) );
  d_ff \prgm_register/genblk1[809].single_DFF  ( .d(
        \prgm_register/or_signal [809]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[809]) );
  d_ff \prgm_register/genblk1[808].single_DFF  ( .d(
        \prgm_register/or_signal [808]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[808]) );
  d_ff \prgm_register/genblk1[807].single_DFF  ( .d(
        \prgm_register/or_signal [807]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[807]) );
  d_ff \prgm_register/genblk1[806].single_DFF  ( .d(
        \prgm_register/or_signal [806]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[806]) );
  d_ff \prgm_register/genblk1[805].single_DFF  ( .d(
        \prgm_register/or_signal [805]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[805]) );
  d_ff \prgm_register/genblk1[804].single_DFF  ( .d(
        \prgm_register/or_signal [804]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[804]) );
  d_ff \prgm_register/genblk1[803].single_DFF  ( .d(
        \prgm_register/or_signal [803]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[803]) );
  d_ff \prgm_register/genblk1[802].single_DFF  ( .d(
        \prgm_register/or_signal [802]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[802]) );
  d_ff \prgm_register/genblk1[801].single_DFF  ( .d(
        \prgm_register/or_signal [801]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[801]) );
  d_ff \prgm_register/genblk1[800].single_DFF  ( .d(
        \prgm_register/or_signal [800]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[800]) );
  d_ff \prgm_register/genblk1[799].single_DFF  ( .d(
        \prgm_register/or_signal [799]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[799]) );
  d_ff \prgm_register/genblk1[798].single_DFF  ( .d(
        \prgm_register/or_signal [798]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[798]) );
  d_ff \prgm_register/genblk1[797].single_DFF  ( .d(
        \prgm_register/or_signal [797]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[797]) );
  d_ff \prgm_register/genblk1[796].single_DFF  ( .d(
        \prgm_register/or_signal [796]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[796]) );
  d_ff \prgm_register/genblk1[795].single_DFF  ( .d(
        \prgm_register/or_signal [795]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[795]) );
  d_ff \prgm_register/genblk1[794].single_DFF  ( .d(
        \prgm_register/or_signal [794]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[794]) );
  d_ff \prgm_register/genblk1[793].single_DFF  ( .d(
        \prgm_register/or_signal [793]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[793]) );
  d_ff \prgm_register/genblk1[792].single_DFF  ( .d(
        \prgm_register/or_signal [792]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[792]) );
  d_ff \prgm_register/genblk1[791].single_DFF  ( .d(
        \prgm_register/or_signal [791]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[791]) );
  d_ff \prgm_register/genblk1[790].single_DFF  ( .d(
        \prgm_register/or_signal [790]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[790]) );
  d_ff \prgm_register/genblk1[789].single_DFF  ( .d(
        \prgm_register/or_signal [789]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[789]) );
  d_ff \prgm_register/genblk1[788].single_DFF  ( .d(
        \prgm_register/or_signal [788]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[788]) );
  d_ff \prgm_register/genblk1[787].single_DFF  ( .d(
        \prgm_register/or_signal [787]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[787]) );
  d_ff \prgm_register/genblk1[786].single_DFF  ( .d(
        \prgm_register/or_signal [786]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[786]) );
  d_ff \prgm_register/genblk1[785].single_DFF  ( .d(
        \prgm_register/or_signal [785]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[785]) );
  d_ff \prgm_register/genblk1[784].single_DFF  ( .d(
        \prgm_register/or_signal [784]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[784]) );
  d_ff \prgm_register/genblk1[783].single_DFF  ( .d(
        \prgm_register/or_signal [783]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[783]) );
  d_ff \prgm_register/genblk1[782].single_DFF  ( .d(
        \prgm_register/or_signal [782]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[782]) );
  d_ff \prgm_register/genblk1[781].single_DFF  ( .d(
        \prgm_register/or_signal [781]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[781]) );
  d_ff \prgm_register/genblk1[780].single_DFF  ( .d(
        \prgm_register/or_signal [780]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[780]) );
  d_ff \prgm_register/genblk1[779].single_DFF  ( .d(
        \prgm_register/or_signal [779]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[779]) );
  d_ff \prgm_register/genblk1[778].single_DFF  ( .d(
        \prgm_register/or_signal [778]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[778]) );
  d_ff \prgm_register/genblk1[777].single_DFF  ( .d(
        \prgm_register/or_signal [777]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[777]) );
  d_ff \prgm_register/genblk1[776].single_DFF  ( .d(
        \prgm_register/or_signal [776]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[776]) );
  d_ff \prgm_register/genblk1[775].single_DFF  ( .d(
        \prgm_register/or_signal [775]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[775]) );
  d_ff \prgm_register/genblk1[774].single_DFF  ( .d(
        \prgm_register/or_signal [774]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[774]) );
  d_ff \prgm_register/genblk1[773].single_DFF  ( .d(
        \prgm_register/or_signal [773]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[773]) );
  d_ff \prgm_register/genblk1[772].single_DFF  ( .d(
        \prgm_register/or_signal [772]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[772]) );
  d_ff \prgm_register/genblk1[771].single_DFF  ( .d(
        \prgm_register/or_signal [771]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[771]) );
  d_ff \prgm_register/genblk1[770].single_DFF  ( .d(
        \prgm_register/or_signal [770]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[770]) );
  d_ff \prgm_register/genblk1[769].single_DFF  ( .d(
        \prgm_register/or_signal [769]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[769]) );
  d_ff \prgm_register/genblk1[768].single_DFF  ( .d(
        \prgm_register/or_signal [768]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[768]) );
  d_ff \prgm_register/genblk1[767].single_DFF  ( .d(
        \prgm_register/or_signal [767]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[767]) );
  d_ff \prgm_register/genblk1[766].single_DFF  ( .d(
        \prgm_register/or_signal [766]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[766]) );
  d_ff \prgm_register/genblk1[765].single_DFF  ( .d(
        \prgm_register/or_signal [765]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[765]) );
  d_ff \prgm_register/genblk1[764].single_DFF  ( .d(
        \prgm_register/or_signal [764]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[764]) );
  d_ff \prgm_register/genblk1[763].single_DFF  ( .d(
        \prgm_register/or_signal [763]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[763]) );
  d_ff \prgm_register/genblk1[762].single_DFF  ( .d(
        \prgm_register/or_signal [762]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[762]) );
  d_ff \prgm_register/genblk1[761].single_DFF  ( .d(
        \prgm_register/or_signal [761]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[761]) );
  d_ff \prgm_register/genblk1[760].single_DFF  ( .d(
        \prgm_register/or_signal [760]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[760]) );
  d_ff \prgm_register/genblk1[759].single_DFF  ( .d(
        \prgm_register/or_signal [759]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[759]) );
  d_ff \prgm_register/genblk1[758].single_DFF  ( .d(
        \prgm_register/or_signal [758]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[758]) );
  d_ff \prgm_register/genblk1[757].single_DFF  ( .d(
        \prgm_register/or_signal [757]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[757]) );
  d_ff \prgm_register/genblk1[756].single_DFF  ( .d(
        \prgm_register/or_signal [756]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[756]) );
  d_ff \prgm_register/genblk1[755].single_DFF  ( .d(
        \prgm_register/or_signal [755]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[755]) );
  d_ff \prgm_register/genblk1[754].single_DFF  ( .d(
        \prgm_register/or_signal [754]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[754]) );
  d_ff \prgm_register/genblk1[753].single_DFF  ( .d(
        \prgm_register/or_signal [753]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[753]) );
  d_ff \prgm_register/genblk1[752].single_DFF  ( .d(
        \prgm_register/or_signal [752]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[752]) );
  d_ff \prgm_register/genblk1[751].single_DFF  ( .d(
        \prgm_register/or_signal [751]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[751]) );
  d_ff \prgm_register/genblk1[750].single_DFF  ( .d(
        \prgm_register/or_signal [750]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[750]) );
  d_ff \prgm_register/genblk1[749].single_DFF  ( .d(
        \prgm_register/or_signal [749]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[749]) );
  d_ff \prgm_register/genblk1[748].single_DFF  ( .d(
        \prgm_register/or_signal [748]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[748]) );
  d_ff \prgm_register/genblk1[747].single_DFF  ( .d(
        \prgm_register/or_signal [747]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[747]) );
  d_ff \prgm_register/genblk1[746].single_DFF  ( .d(
        \prgm_register/or_signal [746]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[746]) );
  d_ff \prgm_register/genblk1[745].single_DFF  ( .d(
        \prgm_register/or_signal [745]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[745]) );
  d_ff \prgm_register/genblk1[744].single_DFF  ( .d(
        \prgm_register/or_signal [744]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[744]) );
  d_ff \prgm_register/genblk1[743].single_DFF  ( .d(
        \prgm_register/or_signal [743]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[743]) );
  d_ff \prgm_register/genblk1[742].single_DFF  ( .d(
        \prgm_register/or_signal [742]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[742]) );
  d_ff \prgm_register/genblk1[741].single_DFF  ( .d(
        \prgm_register/or_signal [741]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[741]) );
  d_ff \prgm_register/genblk1[740].single_DFF  ( .d(
        \prgm_register/or_signal [740]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[740]) );
  d_ff \prgm_register/genblk1[739].single_DFF  ( .d(
        \prgm_register/or_signal [739]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[739]) );
  d_ff \prgm_register/genblk1[738].single_DFF  ( .d(
        \prgm_register/or_signal [738]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[738]) );
  d_ff \prgm_register/genblk1[737].single_DFF  ( .d(
        \prgm_register/or_signal [737]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[737]) );
  d_ff \prgm_register/genblk1[736].single_DFF  ( .d(
        \prgm_register/or_signal [736]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[736]) );
  d_ff \prgm_register/genblk1[735].single_DFF  ( .d(
        \prgm_register/or_signal [735]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[735]) );
  d_ff \prgm_register/genblk1[734].single_DFF  ( .d(
        \prgm_register/or_signal [734]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[734]) );
  d_ff \prgm_register/genblk1[733].single_DFF  ( .d(
        \prgm_register/or_signal [733]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[733]) );
  d_ff \prgm_register/genblk1[732].single_DFF  ( .d(
        \prgm_register/or_signal [732]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[732]) );
  d_ff \prgm_register/genblk1[731].single_DFF  ( .d(
        \prgm_register/or_signal [731]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[731]) );
  d_ff \prgm_register/genblk1[730].single_DFF  ( .d(
        \prgm_register/or_signal [730]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[730]) );
  d_ff \prgm_register/genblk1[729].single_DFF  ( .d(
        \prgm_register/or_signal [729]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[729]) );
  d_ff \prgm_register/genblk1[728].single_DFF  ( .d(
        \prgm_register/or_signal [728]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[728]) );
  d_ff \prgm_register/genblk1[727].single_DFF  ( .d(
        \prgm_register/or_signal [727]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[727]) );
  d_ff \prgm_register/genblk1[726].single_DFF  ( .d(
        \prgm_register/or_signal [726]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[726]) );
  d_ff \prgm_register/genblk1[725].single_DFF  ( .d(
        \prgm_register/or_signal [725]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[725]) );
  d_ff \prgm_register/genblk1[724].single_DFF  ( .d(
        \prgm_register/or_signal [724]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[724]) );
  d_ff \prgm_register/genblk1[723].single_DFF  ( .d(
        \prgm_register/or_signal [723]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[723]) );
  d_ff \prgm_register/genblk1[722].single_DFF  ( .d(
        \prgm_register/or_signal [722]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[722]) );
  d_ff \prgm_register/genblk1[721].single_DFF  ( .d(
        \prgm_register/or_signal [721]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[721]) );
  d_ff \prgm_register/genblk1[720].single_DFF  ( .d(
        \prgm_register/or_signal [720]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[720]) );
  d_ff \prgm_register/genblk1[719].single_DFF  ( .d(
        \prgm_register/or_signal [719]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[719]) );
  d_ff \prgm_register/genblk1[718].single_DFF  ( .d(
        \prgm_register/or_signal [718]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[718]) );
  d_ff \prgm_register/genblk1[717].single_DFF  ( .d(
        \prgm_register/or_signal [717]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[717]) );
  d_ff \prgm_register/genblk1[716].single_DFF  ( .d(
        \prgm_register/or_signal [716]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[716]) );
  d_ff \prgm_register/genblk1[715].single_DFF  ( .d(
        \prgm_register/or_signal [715]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[715]) );
  d_ff \prgm_register/genblk1[714].single_DFF  ( .d(
        \prgm_register/or_signal [714]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[714]) );
  d_ff \prgm_register/genblk1[713].single_DFF  ( .d(
        \prgm_register/or_signal [713]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[713]) );
  d_ff \prgm_register/genblk1[712].single_DFF  ( .d(
        \prgm_register/or_signal [712]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[712]) );
  d_ff \prgm_register/genblk1[711].single_DFF  ( .d(
        \prgm_register/or_signal [711]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[711]) );
  d_ff \prgm_register/genblk1[710].single_DFF  ( .d(
        \prgm_register/or_signal [710]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[710]) );
  d_ff \prgm_register/genblk1[709].single_DFF  ( .d(
        \prgm_register/or_signal [709]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[709]) );
  d_ff \prgm_register/genblk1[708].single_DFF  ( .d(
        \prgm_register/or_signal [708]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[708]) );
  d_ff \prgm_register/genblk1[707].single_DFF  ( .d(
        \prgm_register/or_signal [707]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[707]) );
  d_ff \prgm_register/genblk1[706].single_DFF  ( .d(
        \prgm_register/or_signal [706]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[706]) );
  d_ff \prgm_register/genblk1[705].single_DFF  ( .d(
        \prgm_register/or_signal [705]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[705]) );
  d_ff \prgm_register/genblk1[704].single_DFF  ( .d(
        \prgm_register/or_signal [704]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[704]) );
  d_ff \prgm_register/genblk1[703].single_DFF  ( .d(
        \prgm_register/or_signal [703]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[703]) );
  d_ff \prgm_register/genblk1[702].single_DFF  ( .d(
        \prgm_register/or_signal [702]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[702]) );
  d_ff \prgm_register/genblk1[701].single_DFF  ( .d(
        \prgm_register/or_signal [701]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[701]) );
  d_ff \prgm_register/genblk1[700].single_DFF  ( .d(
        \prgm_register/or_signal [700]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[700]) );
  d_ff \prgm_register/genblk1[699].single_DFF  ( .d(
        \prgm_register/or_signal [699]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[699]) );
  d_ff \prgm_register/genblk1[698].single_DFF  ( .d(
        \prgm_register/or_signal [698]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[698]) );
  d_ff \prgm_register/genblk1[697].single_DFF  ( .d(
        \prgm_register/or_signal [697]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[697]) );
  d_ff \prgm_register/genblk1[696].single_DFF  ( .d(
        \prgm_register/or_signal [696]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[696]) );
  d_ff \prgm_register/genblk1[695].single_DFF  ( .d(
        \prgm_register/or_signal [695]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[695]) );
  d_ff \prgm_register/genblk1[694].single_DFF  ( .d(
        \prgm_register/or_signal [694]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[694]) );
  d_ff \prgm_register/genblk1[693].single_DFF  ( .d(
        \prgm_register/or_signal [693]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[693]) );
  d_ff \prgm_register/genblk1[692].single_DFF  ( .d(
        \prgm_register/or_signal [692]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[692]) );
  d_ff \prgm_register/genblk1[691].single_DFF  ( .d(
        \prgm_register/or_signal [691]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[691]) );
  d_ff \prgm_register/genblk1[690].single_DFF  ( .d(
        \prgm_register/or_signal [690]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[690]) );
  d_ff \prgm_register/genblk1[689].single_DFF  ( .d(
        \prgm_register/or_signal [689]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[689]) );
  d_ff \prgm_register/genblk1[688].single_DFF  ( .d(
        \prgm_register/or_signal [688]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[688]) );
  d_ff \prgm_register/genblk1[687].single_DFF  ( .d(
        \prgm_register/or_signal [687]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[687]) );
  d_ff \prgm_register/genblk1[686].single_DFF  ( .d(
        \prgm_register/or_signal [686]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[686]) );
  d_ff \prgm_register/genblk1[685].single_DFF  ( .d(
        \prgm_register/or_signal [685]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[685]) );
  d_ff \prgm_register/genblk1[684].single_DFF  ( .d(
        \prgm_register/or_signal [684]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[684]) );
  d_ff \prgm_register/genblk1[683].single_DFF  ( .d(
        \prgm_register/or_signal [683]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[683]) );
  d_ff \prgm_register/genblk1[682].single_DFF  ( .d(
        \prgm_register/or_signal [682]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[682]) );
  d_ff \prgm_register/genblk1[681].single_DFF  ( .d(
        \prgm_register/or_signal [681]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[681]) );
  d_ff \prgm_register/genblk1[680].single_DFF  ( .d(
        \prgm_register/or_signal [680]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[680]) );
  d_ff \prgm_register/genblk1[679].single_DFF  ( .d(
        \prgm_register/or_signal [679]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[679]) );
  d_ff \prgm_register/genblk1[678].single_DFF  ( .d(
        \prgm_register/or_signal [678]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[678]) );
  d_ff \prgm_register/genblk1[677].single_DFF  ( .d(
        \prgm_register/or_signal [677]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[677]) );
  d_ff \prgm_register/genblk1[676].single_DFF  ( .d(
        \prgm_register/or_signal [676]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[676]) );
  d_ff \prgm_register/genblk1[675].single_DFF  ( .d(
        \prgm_register/or_signal [675]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[675]) );
  d_ff \prgm_register/genblk1[674].single_DFF  ( .d(
        \prgm_register/or_signal [674]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[674]) );
  d_ff \prgm_register/genblk1[673].single_DFF  ( .d(
        \prgm_register/or_signal [673]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[673]) );
  d_ff \prgm_register/genblk1[672].single_DFF  ( .d(
        \prgm_register/or_signal [672]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[672]) );
  d_ff \prgm_register/genblk1[671].single_DFF  ( .d(
        \prgm_register/or_signal [671]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[671]) );
  d_ff \prgm_register/genblk1[670].single_DFF  ( .d(
        \prgm_register/or_signal [670]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[670]) );
  d_ff \prgm_register/genblk1[669].single_DFF  ( .d(
        \prgm_register/or_signal [669]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[669]) );
  d_ff \prgm_register/genblk1[668].single_DFF  ( .d(
        \prgm_register/or_signal [668]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[668]) );
  d_ff \prgm_register/genblk1[667].single_DFF  ( .d(
        \prgm_register/or_signal [667]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[667]) );
  d_ff \prgm_register/genblk1[666].single_DFF  ( .d(
        \prgm_register/or_signal [666]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[666]) );
  d_ff \prgm_register/genblk1[665].single_DFF  ( .d(
        \prgm_register/or_signal [665]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[665]) );
  d_ff \prgm_register/genblk1[664].single_DFF  ( .d(
        \prgm_register/or_signal [664]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[664]) );
  d_ff \prgm_register/genblk1[663].single_DFF  ( .d(
        \prgm_register/or_signal [663]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[663]) );
  d_ff \prgm_register/genblk1[662].single_DFF  ( .d(
        \prgm_register/or_signal [662]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[662]) );
  d_ff \prgm_register/genblk1[661].single_DFF  ( .d(
        \prgm_register/or_signal [661]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[661]) );
  d_ff \prgm_register/genblk1[660].single_DFF  ( .d(
        \prgm_register/or_signal [660]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[660]) );
  d_ff \prgm_register/genblk1[659].single_DFF  ( .d(
        \prgm_register/or_signal [659]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[659]) );
  d_ff \prgm_register/genblk1[658].single_DFF  ( .d(
        \prgm_register/or_signal [658]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[658]) );
  d_ff \prgm_register/genblk1[657].single_DFF  ( .d(
        \prgm_register/or_signal [657]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[657]) );
  d_ff \prgm_register/genblk1[656].single_DFF  ( .d(
        \prgm_register/or_signal [656]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[656]) );
  d_ff \prgm_register/genblk1[655].single_DFF  ( .d(
        \prgm_register/or_signal [655]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[655]) );
  d_ff \prgm_register/genblk1[654].single_DFF  ( .d(
        \prgm_register/or_signal [654]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[654]) );
  d_ff \prgm_register/genblk1[653].single_DFF  ( .d(
        \prgm_register/or_signal [653]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[653]) );
  d_ff \prgm_register/genblk1[652].single_DFF  ( .d(
        \prgm_register/or_signal [652]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[652]) );
  d_ff \prgm_register/genblk1[651].single_DFF  ( .d(
        \prgm_register/or_signal [651]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[651]) );
  d_ff \prgm_register/genblk1[650].single_DFF  ( .d(
        \prgm_register/or_signal [650]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[650]) );
  d_ff \prgm_register/genblk1[649].single_DFF  ( .d(
        \prgm_register/or_signal [649]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[649]) );
  d_ff \prgm_register/genblk1[648].single_DFF  ( .d(
        \prgm_register/or_signal [648]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[648]) );
  d_ff \prgm_register/genblk1[647].single_DFF  ( .d(
        \prgm_register/or_signal [647]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[647]) );
  d_ff \prgm_register/genblk1[646].single_DFF  ( .d(
        \prgm_register/or_signal [646]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[646]) );
  d_ff \prgm_register/genblk1[645].single_DFF  ( .d(
        \prgm_register/or_signal [645]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[645]) );
  d_ff \prgm_register/genblk1[644].single_DFF  ( .d(
        \prgm_register/or_signal [644]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[644]) );
  d_ff \prgm_register/genblk1[643].single_DFF  ( .d(
        \prgm_register/or_signal [643]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[643]) );
  d_ff \prgm_register/genblk1[642].single_DFF  ( .d(
        \prgm_register/or_signal [642]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[642]) );
  d_ff \prgm_register/genblk1[641].single_DFF  ( .d(
        \prgm_register/or_signal [641]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[641]) );
  d_ff \prgm_register/genblk1[640].single_DFF  ( .d(
        \prgm_register/or_signal [640]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[640]) );
  d_ff \prgm_register/genblk1[639].single_DFF  ( .d(
        \prgm_register/or_signal [639]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[639]) );
  d_ff \prgm_register/genblk1[638].single_DFF  ( .d(
        \prgm_register/or_signal [638]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[638]) );
  d_ff \prgm_register/genblk1[637].single_DFF  ( .d(
        \prgm_register/or_signal [637]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[637]) );
  d_ff \prgm_register/genblk1[636].single_DFF  ( .d(
        \prgm_register/or_signal [636]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[636]) );
  d_ff \prgm_register/genblk1[635].single_DFF  ( .d(
        \prgm_register/or_signal [635]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[635]) );
  d_ff \prgm_register/genblk1[634].single_DFF  ( .d(
        \prgm_register/or_signal [634]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[634]) );
  d_ff \prgm_register/genblk1[633].single_DFF  ( .d(
        \prgm_register/or_signal [633]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[633]) );
  d_ff \prgm_register/genblk1[632].single_DFF  ( .d(
        \prgm_register/or_signal [632]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[632]) );
  d_ff \prgm_register/genblk1[631].single_DFF  ( .d(
        \prgm_register/or_signal [631]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[631]) );
  d_ff \prgm_register/genblk1[630].single_DFF  ( .d(
        \prgm_register/or_signal [630]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[630]) );
  d_ff \prgm_register/genblk1[629].single_DFF  ( .d(
        \prgm_register/or_signal [629]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[629]) );
  d_ff \prgm_register/genblk1[628].single_DFF  ( .d(
        \prgm_register/or_signal [628]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[628]) );
  d_ff \prgm_register/genblk1[627].single_DFF  ( .d(
        \prgm_register/or_signal [627]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[627]) );
  d_ff \prgm_register/genblk1[626].single_DFF  ( .d(
        \prgm_register/or_signal [626]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[626]) );
  d_ff \prgm_register/genblk1[625].single_DFF  ( .d(
        \prgm_register/or_signal [625]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[625]) );
  d_ff \prgm_register/genblk1[624].single_DFF  ( .d(
        \prgm_register/or_signal [624]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[624]) );
  d_ff \prgm_register/genblk1[623].single_DFF  ( .d(
        \prgm_register/or_signal [623]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[623]) );
  d_ff \prgm_register/genblk1[622].single_DFF  ( .d(
        \prgm_register/or_signal [622]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[622]) );
  d_ff \prgm_register/genblk1[621].single_DFF  ( .d(
        \prgm_register/or_signal [621]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[621]) );
  d_ff \prgm_register/genblk1[620].single_DFF  ( .d(
        \prgm_register/or_signal [620]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[620]) );
  d_ff \prgm_register/genblk1[619].single_DFF  ( .d(
        \prgm_register/or_signal [619]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[619]) );
  d_ff \prgm_register/genblk1[618].single_DFF  ( .d(
        \prgm_register/or_signal [618]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[618]) );
  d_ff \prgm_register/genblk1[617].single_DFF  ( .d(
        \prgm_register/or_signal [617]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[617]) );
  d_ff \prgm_register/genblk1[616].single_DFF  ( .d(
        \prgm_register/or_signal [616]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[616]) );
  d_ff \prgm_register/genblk1[615].single_DFF  ( .d(
        \prgm_register/or_signal [615]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[615]) );
  d_ff \prgm_register/genblk1[614].single_DFF  ( .d(
        \prgm_register/or_signal [614]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[614]) );
  d_ff \prgm_register/genblk1[613].single_DFF  ( .d(
        \prgm_register/or_signal [613]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[613]) );
  d_ff \prgm_register/genblk1[612].single_DFF  ( .d(
        \prgm_register/or_signal [612]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[612]) );
  d_ff \prgm_register/genblk1[611].single_DFF  ( .d(
        \prgm_register/or_signal [611]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[611]) );
  d_ff \prgm_register/genblk1[610].single_DFF  ( .d(
        \prgm_register/or_signal [610]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[610]) );
  d_ff \prgm_register/genblk1[609].single_DFF  ( .d(
        \prgm_register/or_signal [609]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[609]) );
  d_ff \prgm_register/genblk1[608].single_DFF  ( .d(
        \prgm_register/or_signal [608]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[608]) );
  d_ff \prgm_register/genblk1[607].single_DFF  ( .d(
        \prgm_register/or_signal [607]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[607]) );
  d_ff \prgm_register/genblk1[606].single_DFF  ( .d(
        \prgm_register/or_signal [606]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[606]) );
  d_ff \prgm_register/genblk1[605].single_DFF  ( .d(
        \prgm_register/or_signal [605]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[605]) );
  d_ff \prgm_register/genblk1[604].single_DFF  ( .d(
        \prgm_register/or_signal [604]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[604]) );
  d_ff \prgm_register/genblk1[603].single_DFF  ( .d(
        \prgm_register/or_signal [603]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[603]) );
  d_ff \prgm_register/genblk1[602].single_DFF  ( .d(
        \prgm_register/or_signal [602]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[602]) );
  d_ff \prgm_register/genblk1[601].single_DFF  ( .d(
        \prgm_register/or_signal [601]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[601]) );
  d_ff \prgm_register/genblk1[600].single_DFF  ( .d(
        \prgm_register/or_signal [600]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[600]) );
  d_ff \prgm_register/genblk1[599].single_DFF  ( .d(
        \prgm_register/or_signal [599]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[599]) );
  d_ff \prgm_register/genblk1[598].single_DFF  ( .d(
        \prgm_register/or_signal [598]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[598]) );
  d_ff \prgm_register/genblk1[597].single_DFF  ( .d(
        \prgm_register/or_signal [597]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[597]) );
  d_ff \prgm_register/genblk1[596].single_DFF  ( .d(
        \prgm_register/or_signal [596]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[596]) );
  d_ff \prgm_register/genblk1[595].single_DFF  ( .d(
        \prgm_register/or_signal [595]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[595]) );
  d_ff \prgm_register/genblk1[594].single_DFF  ( .d(
        \prgm_register/or_signal [594]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[594]) );
  d_ff \prgm_register/genblk1[593].single_DFF  ( .d(
        \prgm_register/or_signal [593]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[593]) );
  d_ff \prgm_register/genblk1[592].single_DFF  ( .d(
        \prgm_register/or_signal [592]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[592]) );
  d_ff \prgm_register/genblk1[591].single_DFF  ( .d(
        \prgm_register/or_signal [591]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[591]) );
  d_ff \prgm_register/genblk1[590].single_DFF  ( .d(
        \prgm_register/or_signal [590]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[590]) );
  d_ff \prgm_register/genblk1[589].single_DFF  ( .d(
        \prgm_register/or_signal [589]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[589]) );
  d_ff \prgm_register/genblk1[588].single_DFF  ( .d(
        \prgm_register/or_signal [588]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[588]) );
  d_ff \prgm_register/genblk1[587].single_DFF  ( .d(
        \prgm_register/or_signal [587]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[587]) );
  d_ff \prgm_register/genblk1[586].single_DFF  ( .d(
        \prgm_register/or_signal [586]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[586]) );
  d_ff \prgm_register/genblk1[585].single_DFF  ( .d(
        \prgm_register/or_signal [585]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[585]) );
  d_ff \prgm_register/genblk1[584].single_DFF  ( .d(
        \prgm_register/or_signal [584]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[584]) );
  d_ff \prgm_register/genblk1[583].single_DFF  ( .d(
        \prgm_register/or_signal [583]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[583]) );
  d_ff \prgm_register/genblk1[582].single_DFF  ( .d(
        \prgm_register/or_signal [582]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[582]) );
  d_ff \prgm_register/genblk1[581].single_DFF  ( .d(
        \prgm_register/or_signal [581]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[581]) );
  d_ff \prgm_register/genblk1[580].single_DFF  ( .d(
        \prgm_register/or_signal [580]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[580]) );
  d_ff \prgm_register/genblk1[579].single_DFF  ( .d(
        \prgm_register/or_signal [579]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[579]) );
  d_ff \prgm_register/genblk1[578].single_DFF  ( .d(
        \prgm_register/or_signal [578]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[578]) );
  d_ff \prgm_register/genblk1[577].single_DFF  ( .d(
        \prgm_register/or_signal [577]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[577]) );
  d_ff \prgm_register/genblk1[576].single_DFF  ( .d(
        \prgm_register/or_signal [576]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[576]) );
  d_ff \prgm_register/genblk1[575].single_DFF  ( .d(
        \prgm_register/or_signal [575]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[575]) );
  d_ff \prgm_register/genblk1[574].single_DFF  ( .d(
        \prgm_register/or_signal [574]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[574]) );
  d_ff \prgm_register/genblk1[573].single_DFF  ( .d(
        \prgm_register/or_signal [573]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[573]) );
  d_ff \prgm_register/genblk1[572].single_DFF  ( .d(
        \prgm_register/or_signal [572]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[572]) );
  d_ff \prgm_register/genblk1[571].single_DFF  ( .d(
        \prgm_register/or_signal [571]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[571]) );
  d_ff \prgm_register/genblk1[570].single_DFF  ( .d(
        \prgm_register/or_signal [570]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[570]) );
  d_ff \prgm_register/genblk1[569].single_DFF  ( .d(
        \prgm_register/or_signal [569]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[569]) );
  d_ff \prgm_register/genblk1[568].single_DFF  ( .d(
        \prgm_register/or_signal [568]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[568]) );
  d_ff \prgm_register/genblk1[567].single_DFF  ( .d(
        \prgm_register/or_signal [567]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[567]) );
  d_ff \prgm_register/genblk1[566].single_DFF  ( .d(
        \prgm_register/or_signal [566]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[566]) );
  d_ff \prgm_register/genblk1[565].single_DFF  ( .d(
        \prgm_register/or_signal [565]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[565]) );
  d_ff \prgm_register/genblk1[564].single_DFF  ( .d(
        \prgm_register/or_signal [564]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[564]) );
  d_ff \prgm_register/genblk1[563].single_DFF  ( .d(
        \prgm_register/or_signal [563]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[563]) );
  d_ff \prgm_register/genblk1[562].single_DFF  ( .d(
        \prgm_register/or_signal [562]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[562]) );
  d_ff \prgm_register/genblk1[561].single_DFF  ( .d(
        \prgm_register/or_signal [561]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[561]) );
  d_ff \prgm_register/genblk1[560].single_DFF  ( .d(
        \prgm_register/or_signal [560]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[560]) );
  d_ff \prgm_register/genblk1[559].single_DFF  ( .d(
        \prgm_register/or_signal [559]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[559]) );
  d_ff \prgm_register/genblk1[558].single_DFF  ( .d(
        \prgm_register/or_signal [558]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[558]) );
  d_ff \prgm_register/genblk1[557].single_DFF  ( .d(
        \prgm_register/or_signal [557]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[557]) );
  d_ff \prgm_register/genblk1[556].single_DFF  ( .d(
        \prgm_register/or_signal [556]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[556]) );
  d_ff \prgm_register/genblk1[555].single_DFF  ( .d(
        \prgm_register/or_signal [555]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[555]) );
  d_ff \prgm_register/genblk1[554].single_DFF  ( .d(
        \prgm_register/or_signal [554]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[554]) );
  d_ff \prgm_register/genblk1[553].single_DFF  ( .d(
        \prgm_register/or_signal [553]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[553]) );
  d_ff \prgm_register/genblk1[552].single_DFF  ( .d(
        \prgm_register/or_signal [552]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[552]) );
  d_ff \prgm_register/genblk1[551].single_DFF  ( .d(
        \prgm_register/or_signal [551]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[551]) );
  d_ff \prgm_register/genblk1[550].single_DFF  ( .d(
        \prgm_register/or_signal [550]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[550]) );
  d_ff \prgm_register/genblk1[549].single_DFF  ( .d(
        \prgm_register/or_signal [549]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[549]) );
  d_ff \prgm_register/genblk1[548].single_DFF  ( .d(
        \prgm_register/or_signal [548]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[548]) );
  d_ff \prgm_register/genblk1[547].single_DFF  ( .d(
        \prgm_register/or_signal [547]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[547]) );
  d_ff \prgm_register/genblk1[546].single_DFF  ( .d(
        \prgm_register/or_signal [546]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[546]) );
  d_ff \prgm_register/genblk1[545].single_DFF  ( .d(
        \prgm_register/or_signal [545]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[545]) );
  d_ff \prgm_register/genblk1[544].single_DFF  ( .d(
        \prgm_register/or_signal [544]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[544]) );
  d_ff \prgm_register/genblk1[543].single_DFF  ( .d(
        \prgm_register/or_signal [543]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[543]) );
  d_ff \prgm_register/genblk1[542].single_DFF  ( .d(
        \prgm_register/or_signal [542]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[542]) );
  d_ff \prgm_register/genblk1[541].single_DFF  ( .d(
        \prgm_register/or_signal [541]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[541]) );
  d_ff \prgm_register/genblk1[540].single_DFF  ( .d(
        \prgm_register/or_signal [540]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[540]) );
  d_ff \prgm_register/genblk1[539].single_DFF  ( .d(
        \prgm_register/or_signal [539]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[539]) );
  d_ff \prgm_register/genblk1[538].single_DFF  ( .d(
        \prgm_register/or_signal [538]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[538]) );
  d_ff \prgm_register/genblk1[537].single_DFF  ( .d(
        \prgm_register/or_signal [537]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[537]) );
  d_ff \prgm_register/genblk1[536].single_DFF  ( .d(
        \prgm_register/or_signal [536]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[536]) );
  d_ff \prgm_register/genblk1[535].single_DFF  ( .d(
        \prgm_register/or_signal [535]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[535]) );
  d_ff \prgm_register/genblk1[534].single_DFF  ( .d(
        \prgm_register/or_signal [534]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[534]) );
  d_ff \prgm_register/genblk1[533].single_DFF  ( .d(
        \prgm_register/or_signal [533]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[533]) );
  d_ff \prgm_register/genblk1[532].single_DFF  ( .d(
        \prgm_register/or_signal [532]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[532]) );
  d_ff \prgm_register/genblk1[531].single_DFF  ( .d(
        \prgm_register/or_signal [531]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[531]) );
  d_ff \prgm_register/genblk1[530].single_DFF  ( .d(
        \prgm_register/or_signal [530]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[530]) );
  d_ff \prgm_register/genblk1[529].single_DFF  ( .d(
        \prgm_register/or_signal [529]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[529]) );
  d_ff \prgm_register/genblk1[528].single_DFF  ( .d(
        \prgm_register/or_signal [528]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[528]) );
  d_ff \prgm_register/genblk1[527].single_DFF  ( .d(
        \prgm_register/or_signal [527]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[527]) );
  d_ff \prgm_register/genblk1[526].single_DFF  ( .d(
        \prgm_register/or_signal [526]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[526]) );
  d_ff \prgm_register/genblk1[525].single_DFF  ( .d(
        \prgm_register/or_signal [525]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[525]) );
  d_ff \prgm_register/genblk1[524].single_DFF  ( .d(
        \prgm_register/or_signal [524]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[524]) );
  d_ff \prgm_register/genblk1[523].single_DFF  ( .d(
        \prgm_register/or_signal [523]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[523]) );
  d_ff \prgm_register/genblk1[522].single_DFF  ( .d(
        \prgm_register/or_signal [522]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[522]) );
  d_ff \prgm_register/genblk1[521].single_DFF  ( .d(
        \prgm_register/or_signal [521]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[521]) );
  d_ff \prgm_register/genblk1[520].single_DFF  ( .d(
        \prgm_register/or_signal [520]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[520]) );
  d_ff \prgm_register/genblk1[519].single_DFF  ( .d(
        \prgm_register/or_signal [519]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[519]) );
  d_ff \prgm_register/genblk1[518].single_DFF  ( .d(
        \prgm_register/or_signal [518]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[518]) );
  d_ff \prgm_register/genblk1[517].single_DFF  ( .d(
        \prgm_register/or_signal [517]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[517]) );
  d_ff \prgm_register/genblk1[516].single_DFF  ( .d(
        \prgm_register/or_signal [516]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[516]) );
  d_ff \prgm_register/genblk1[515].single_DFF  ( .d(
        \prgm_register/or_signal [515]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[515]) );
  d_ff \prgm_register/genblk1[514].single_DFF  ( .d(
        \prgm_register/or_signal [514]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[514]) );
  d_ff \prgm_register/genblk1[513].single_DFF  ( .d(
        \prgm_register/or_signal [513]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[513]) );
  d_ff \prgm_register/genblk1[512].single_DFF  ( .d(
        \prgm_register/or_signal [512]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[512]) );
  d_ff \prgm_register/genblk1[511].single_DFF  ( .d(
        \prgm_register/or_signal [511]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[511]) );
  d_ff \prgm_register/genblk1[510].single_DFF  ( .d(
        \prgm_register/or_signal [510]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[510]) );
  d_ff \prgm_register/genblk1[509].single_DFF  ( .d(
        \prgm_register/or_signal [509]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[509]) );
  d_ff \prgm_register/genblk1[508].single_DFF  ( .d(
        \prgm_register/or_signal [508]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[508]) );
  d_ff \prgm_register/genblk1[507].single_DFF  ( .d(
        \prgm_register/or_signal [507]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[507]) );
  d_ff \prgm_register/genblk1[506].single_DFF  ( .d(
        \prgm_register/or_signal [506]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[506]) );
  d_ff \prgm_register/genblk1[505].single_DFF  ( .d(
        \prgm_register/or_signal [505]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[505]) );
  d_ff \prgm_register/genblk1[504].single_DFF  ( .d(
        \prgm_register/or_signal [504]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[504]) );
  d_ff \prgm_register/genblk1[503].single_DFF  ( .d(
        \prgm_register/or_signal [503]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[503]) );
  d_ff \prgm_register/genblk1[502].single_DFF  ( .d(
        \prgm_register/or_signal [502]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[502]) );
  d_ff \prgm_register/genblk1[501].single_DFF  ( .d(
        \prgm_register/or_signal [501]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[501]) );
  d_ff \prgm_register/genblk1[500].single_DFF  ( .d(
        \prgm_register/or_signal [500]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[500]) );
  d_ff \prgm_register/genblk1[499].single_DFF  ( .d(
        \prgm_register/or_signal [499]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[499]) );
  d_ff \prgm_register/genblk1[498].single_DFF  ( .d(
        \prgm_register/or_signal [498]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[498]) );
  d_ff \prgm_register/genblk1[497].single_DFF  ( .d(
        \prgm_register/or_signal [497]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[497]) );
  d_ff \prgm_register/genblk1[496].single_DFF  ( .d(
        \prgm_register/or_signal [496]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[496]) );
  d_ff \prgm_register/genblk1[495].single_DFF  ( .d(
        \prgm_register/or_signal [495]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[495]) );
  d_ff \prgm_register/genblk1[494].single_DFF  ( .d(
        \prgm_register/or_signal [494]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[494]) );
  d_ff \prgm_register/genblk1[493].single_DFF  ( .d(
        \prgm_register/or_signal [493]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[493]) );
  d_ff \prgm_register/genblk1[492].single_DFF  ( .d(
        \prgm_register/or_signal [492]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[492]) );
  d_ff \prgm_register/genblk1[491].single_DFF  ( .d(
        \prgm_register/or_signal [491]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[491]) );
  d_ff \prgm_register/genblk1[490].single_DFF  ( .d(
        \prgm_register/or_signal [490]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[490]) );
  d_ff \prgm_register/genblk1[489].single_DFF  ( .d(
        \prgm_register/or_signal [489]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[489]) );
  d_ff \prgm_register/genblk1[488].single_DFF  ( .d(
        \prgm_register/or_signal [488]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[488]) );
  d_ff \prgm_register/genblk1[487].single_DFF  ( .d(
        \prgm_register/or_signal [487]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[487]) );
  d_ff \prgm_register/genblk1[486].single_DFF  ( .d(
        \prgm_register/or_signal [486]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[486]) );
  d_ff \prgm_register/genblk1[485].single_DFF  ( .d(
        \prgm_register/or_signal [485]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[485]) );
  d_ff \prgm_register/genblk1[484].single_DFF  ( .d(
        \prgm_register/or_signal [484]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[484]) );
  d_ff \prgm_register/genblk1[483].single_DFF  ( .d(
        \prgm_register/or_signal [483]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[483]) );
  d_ff \prgm_register/genblk1[482].single_DFF  ( .d(
        \prgm_register/or_signal [482]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[482]) );
  d_ff \prgm_register/genblk1[481].single_DFF  ( .d(
        \prgm_register/or_signal [481]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[481]) );
  d_ff \prgm_register/genblk1[480].single_DFF  ( .d(
        \prgm_register/or_signal [480]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[480]) );
  d_ff \prgm_register/genblk1[479].single_DFF  ( .d(
        \prgm_register/or_signal [479]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[479]) );
  d_ff \prgm_register/genblk1[478].single_DFF  ( .d(
        \prgm_register/or_signal [478]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[478]) );
  d_ff \prgm_register/genblk1[477].single_DFF  ( .d(
        \prgm_register/or_signal [477]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[477]) );
  d_ff \prgm_register/genblk1[476].single_DFF  ( .d(
        \prgm_register/or_signal [476]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[476]) );
  d_ff \prgm_register/genblk1[475].single_DFF  ( .d(
        \prgm_register/or_signal [475]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[475]) );
  d_ff \prgm_register/genblk1[474].single_DFF  ( .d(
        \prgm_register/or_signal [474]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[474]) );
  d_ff \prgm_register/genblk1[473].single_DFF  ( .d(
        \prgm_register/or_signal [473]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[473]) );
  d_ff \prgm_register/genblk1[472].single_DFF  ( .d(
        \prgm_register/or_signal [472]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[472]) );
  d_ff \prgm_register/genblk1[471].single_DFF  ( .d(
        \prgm_register/or_signal [471]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[471]) );
  d_ff \prgm_register/genblk1[470].single_DFF  ( .d(
        \prgm_register/or_signal [470]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[470]) );
  d_ff \prgm_register/genblk1[469].single_DFF  ( .d(
        \prgm_register/or_signal [469]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[469]) );
  d_ff \prgm_register/genblk1[468].single_DFF  ( .d(
        \prgm_register/or_signal [468]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[468]) );
  d_ff \prgm_register/genblk1[467].single_DFF  ( .d(
        \prgm_register/or_signal [467]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[467]) );
  d_ff \prgm_register/genblk1[466].single_DFF  ( .d(
        \prgm_register/or_signal [466]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[466]) );
  d_ff \prgm_register/genblk1[465].single_DFF  ( .d(
        \prgm_register/or_signal [465]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[465]) );
  d_ff \prgm_register/genblk1[464].single_DFF  ( .d(
        \prgm_register/or_signal [464]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[464]) );
  d_ff \prgm_register/genblk1[463].single_DFF  ( .d(
        \prgm_register/or_signal [463]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[463]) );
  d_ff \prgm_register/genblk1[462].single_DFF  ( .d(
        \prgm_register/or_signal [462]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[462]) );
  d_ff \prgm_register/genblk1[461].single_DFF  ( .d(
        \prgm_register/or_signal [461]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[461]) );
  d_ff \prgm_register/genblk1[460].single_DFF  ( .d(
        \prgm_register/or_signal [460]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[460]) );
  d_ff \prgm_register/genblk1[459].single_DFF  ( .d(
        \prgm_register/or_signal [459]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[459]) );
  d_ff \prgm_register/genblk1[458].single_DFF  ( .d(
        \prgm_register/or_signal [458]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[458]) );
  d_ff \prgm_register/genblk1[457].single_DFF  ( .d(
        \prgm_register/or_signal [457]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[457]) );
  d_ff \prgm_register/genblk1[456].single_DFF  ( .d(
        \prgm_register/or_signal [456]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[456]) );
  d_ff \prgm_register/genblk1[455].single_DFF  ( .d(
        \prgm_register/or_signal [455]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[455]) );
  d_ff \prgm_register/genblk1[454].single_DFF  ( .d(
        \prgm_register/or_signal [454]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[454]) );
  d_ff \prgm_register/genblk1[453].single_DFF  ( .d(
        \prgm_register/or_signal [453]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[453]) );
  d_ff \prgm_register/genblk1[452].single_DFF  ( .d(
        \prgm_register/or_signal [452]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[452]) );
  d_ff \prgm_register/genblk1[451].single_DFF  ( .d(
        \prgm_register/or_signal [451]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[451]) );
  d_ff \prgm_register/genblk1[450].single_DFF  ( .d(
        \prgm_register/or_signal [450]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[450]) );
  d_ff \prgm_register/genblk1[449].single_DFF  ( .d(
        \prgm_register/or_signal [449]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[449]) );
  d_ff \prgm_register/genblk1[448].single_DFF  ( .d(
        \prgm_register/or_signal [448]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[448]) );
  d_ff \prgm_register/genblk1[447].single_DFF  ( .d(
        \prgm_register/or_signal [447]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[447]) );
  d_ff \prgm_register/genblk1[446].single_DFF  ( .d(
        \prgm_register/or_signal [446]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[446]) );
  d_ff \prgm_register/genblk1[445].single_DFF  ( .d(
        \prgm_register/or_signal [445]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[445]) );
  d_ff \prgm_register/genblk1[444].single_DFF  ( .d(
        \prgm_register/or_signal [444]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[444]) );
  d_ff \prgm_register/genblk1[443].single_DFF  ( .d(
        \prgm_register/or_signal [443]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[443]) );
  d_ff \prgm_register/genblk1[442].single_DFF  ( .d(
        \prgm_register/or_signal [442]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[442]) );
  d_ff \prgm_register/genblk1[441].single_DFF  ( .d(
        \prgm_register/or_signal [441]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[441]) );
  d_ff \prgm_register/genblk1[440].single_DFF  ( .d(
        \prgm_register/or_signal [440]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[440]) );
  d_ff \prgm_register/genblk1[439].single_DFF  ( .d(
        \prgm_register/or_signal [439]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[439]) );
  d_ff \prgm_register/genblk1[438].single_DFF  ( .d(
        \prgm_register/or_signal [438]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[438]) );
  d_ff \prgm_register/genblk1[437].single_DFF  ( .d(
        \prgm_register/or_signal [437]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[437]) );
  d_ff \prgm_register/genblk1[436].single_DFF  ( .d(
        \prgm_register/or_signal [436]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[436]) );
  d_ff \prgm_register/genblk1[435].single_DFF  ( .d(
        \prgm_register/or_signal [435]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[435]) );
  d_ff \prgm_register/genblk1[434].single_DFF  ( .d(
        \prgm_register/or_signal [434]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[434]) );
  d_ff \prgm_register/genblk1[433].single_DFF  ( .d(
        \prgm_register/or_signal [433]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[433]) );
  d_ff \prgm_register/genblk1[432].single_DFF  ( .d(
        \prgm_register/or_signal [432]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[432]) );
  d_ff \prgm_register/genblk1[431].single_DFF  ( .d(
        \prgm_register/or_signal [431]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[431]) );
  d_ff \prgm_register/genblk1[430].single_DFF  ( .d(
        \prgm_register/or_signal [430]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[430]) );
  d_ff \prgm_register/genblk1[429].single_DFF  ( .d(
        \prgm_register/or_signal [429]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[429]) );
  d_ff \prgm_register/genblk1[428].single_DFF  ( .d(
        \prgm_register/or_signal [428]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[428]) );
  d_ff \prgm_register/genblk1[427].single_DFF  ( .d(
        \prgm_register/or_signal [427]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[427]) );
  d_ff \prgm_register/genblk1[426].single_DFF  ( .d(
        \prgm_register/or_signal [426]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[426]) );
  d_ff \prgm_register/genblk1[425].single_DFF  ( .d(
        \prgm_register/or_signal [425]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[425]) );
  d_ff \prgm_register/genblk1[424].single_DFF  ( .d(
        \prgm_register/or_signal [424]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[424]) );
  d_ff \prgm_register/genblk1[423].single_DFF  ( .d(
        \prgm_register/or_signal [423]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[423]) );
  d_ff \prgm_register/genblk1[422].single_DFF  ( .d(
        \prgm_register/or_signal [422]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[422]) );
  d_ff \prgm_register/genblk1[421].single_DFF  ( .d(
        \prgm_register/or_signal [421]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[421]) );
  d_ff \prgm_register/genblk1[420].single_DFF  ( .d(
        \prgm_register/or_signal [420]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[420]) );
  d_ff \prgm_register/genblk1[419].single_DFF  ( .d(
        \prgm_register/or_signal [419]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[419]) );
  d_ff \prgm_register/genblk1[418].single_DFF  ( .d(
        \prgm_register/or_signal [418]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[418]) );
  d_ff \prgm_register/genblk1[417].single_DFF  ( .d(
        \prgm_register/or_signal [417]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[417]) );
  d_ff \prgm_register/genblk1[416].single_DFF  ( .d(
        \prgm_register/or_signal [416]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[416]) );
  d_ff \prgm_register/genblk1[415].single_DFF  ( .d(
        \prgm_register/or_signal [415]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[415]) );
  d_ff \prgm_register/genblk1[414].single_DFF  ( .d(
        \prgm_register/or_signal [414]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[414]) );
  d_ff \prgm_register/genblk1[413].single_DFF  ( .d(
        \prgm_register/or_signal [413]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[413]) );
  d_ff \prgm_register/genblk1[412].single_DFF  ( .d(
        \prgm_register/or_signal [412]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[412]) );
  d_ff \prgm_register/genblk1[411].single_DFF  ( .d(
        \prgm_register/or_signal [411]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[411]) );
  d_ff \prgm_register/genblk1[410].single_DFF  ( .d(
        \prgm_register/or_signal [410]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[410]) );
  d_ff \prgm_register/genblk1[409].single_DFF  ( .d(
        \prgm_register/or_signal [409]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[409]) );
  d_ff \prgm_register/genblk1[408].single_DFF  ( .d(
        \prgm_register/or_signal [408]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[408]) );
  d_ff \prgm_register/genblk1[407].single_DFF  ( .d(
        \prgm_register/or_signal [407]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[407]) );
  d_ff \prgm_register/genblk1[406].single_DFF  ( .d(
        \prgm_register/or_signal [406]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[406]) );
  d_ff \prgm_register/genblk1[405].single_DFF  ( .d(
        \prgm_register/or_signal [405]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[405]) );
  d_ff \prgm_register/genblk1[404].single_DFF  ( .d(
        \prgm_register/or_signal [404]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[404]) );
  d_ff \prgm_register/genblk1[403].single_DFF  ( .d(
        \prgm_register/or_signal [403]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[403]) );
  d_ff \prgm_register/genblk1[402].single_DFF  ( .d(
        \prgm_register/or_signal [402]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[402]) );
  d_ff \prgm_register/genblk1[401].single_DFF  ( .d(
        \prgm_register/or_signal [401]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[401]) );
  d_ff \prgm_register/genblk1[400].single_DFF  ( .d(
        \prgm_register/or_signal [400]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[400]) );
  d_ff \prgm_register/genblk1[399].single_DFF  ( .d(
        \prgm_register/or_signal [399]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[399]) );
  d_ff \prgm_register/genblk1[398].single_DFF  ( .d(
        \prgm_register/or_signal [398]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[398]) );
  d_ff \prgm_register/genblk1[397].single_DFF  ( .d(
        \prgm_register/or_signal [397]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[397]) );
  d_ff \prgm_register/genblk1[396].single_DFF  ( .d(
        \prgm_register/or_signal [396]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[396]) );
  d_ff \prgm_register/genblk1[395].single_DFF  ( .d(
        \prgm_register/or_signal [395]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[395]) );
  d_ff \prgm_register/genblk1[394].single_DFF  ( .d(
        \prgm_register/or_signal [394]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[394]) );
  d_ff \prgm_register/genblk1[393].single_DFF  ( .d(
        \prgm_register/or_signal [393]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[393]) );
  d_ff \prgm_register/genblk1[392].single_DFF  ( .d(
        \prgm_register/or_signal [392]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[392]) );
  d_ff \prgm_register/genblk1[391].single_DFF  ( .d(
        \prgm_register/or_signal [391]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[391]) );
  d_ff \prgm_register/genblk1[390].single_DFF  ( .d(
        \prgm_register/or_signal [390]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[390]) );
  d_ff \prgm_register/genblk1[389].single_DFF  ( .d(
        \prgm_register/or_signal [389]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[389]) );
  d_ff \prgm_register/genblk1[388].single_DFF  ( .d(
        \prgm_register/or_signal [388]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[388]) );
  d_ff \prgm_register/genblk1[387].single_DFF  ( .d(
        \prgm_register/or_signal [387]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[387]) );
  d_ff \prgm_register/genblk1[386].single_DFF  ( .d(
        \prgm_register/or_signal [386]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[386]) );
  d_ff \prgm_register/genblk1[385].single_DFF  ( .d(
        \prgm_register/or_signal [385]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[385]) );
  d_ff \prgm_register/genblk1[384].single_DFF  ( .d(
        \prgm_register/or_signal [384]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[384]) );
  d_ff \prgm_register/genblk1[383].single_DFF  ( .d(
        \prgm_register/or_signal [383]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[383]) );
  d_ff \prgm_register/genblk1[382].single_DFF  ( .d(
        \prgm_register/or_signal [382]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[382]) );
  d_ff \prgm_register/genblk1[381].single_DFF  ( .d(
        \prgm_register/or_signal [381]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[381]) );
  d_ff \prgm_register/genblk1[380].single_DFF  ( .d(
        \prgm_register/or_signal [380]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[380]) );
  d_ff \prgm_register/genblk1[379].single_DFF  ( .d(
        \prgm_register/or_signal [379]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[379]) );
  d_ff \prgm_register/genblk1[378].single_DFF  ( .d(
        \prgm_register/or_signal [378]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[378]) );
  d_ff \prgm_register/genblk1[377].single_DFF  ( .d(
        \prgm_register/or_signal [377]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[377]) );
  d_ff \prgm_register/genblk1[376].single_DFF  ( .d(
        \prgm_register/or_signal [376]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[376]) );
  d_ff \prgm_register/genblk1[375].single_DFF  ( .d(
        \prgm_register/or_signal [375]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[375]) );
  d_ff \prgm_register/genblk1[374].single_DFF  ( .d(
        \prgm_register/or_signal [374]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[374]) );
  d_ff \prgm_register/genblk1[373].single_DFF  ( .d(
        \prgm_register/or_signal [373]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[373]) );
  d_ff \prgm_register/genblk1[372].single_DFF  ( .d(
        \prgm_register/or_signal [372]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[372]) );
  d_ff \prgm_register/genblk1[371].single_DFF  ( .d(
        \prgm_register/or_signal [371]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[371]) );
  d_ff \prgm_register/genblk1[370].single_DFF  ( .d(
        \prgm_register/or_signal [370]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[370]) );
  d_ff \prgm_register/genblk1[369].single_DFF  ( .d(
        \prgm_register/or_signal [369]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[369]) );
  d_ff \prgm_register/genblk1[368].single_DFF  ( .d(
        \prgm_register/or_signal [368]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[368]) );
  d_ff \prgm_register/genblk1[367].single_DFF  ( .d(
        \prgm_register/or_signal [367]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[367]) );
  d_ff \prgm_register/genblk1[366].single_DFF  ( .d(
        \prgm_register/or_signal [366]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[366]) );
  d_ff \prgm_register/genblk1[365].single_DFF  ( .d(
        \prgm_register/or_signal [365]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[365]) );
  d_ff \prgm_register/genblk1[364].single_DFF  ( .d(
        \prgm_register/or_signal [364]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[364]) );
  d_ff \prgm_register/genblk1[363].single_DFF  ( .d(
        \prgm_register/or_signal [363]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[363]) );
  d_ff \prgm_register/genblk1[362].single_DFF  ( .d(
        \prgm_register/or_signal [362]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[362]) );
  d_ff \prgm_register/genblk1[361].single_DFF  ( .d(
        \prgm_register/or_signal [361]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[361]) );
  d_ff \prgm_register/genblk1[360].single_DFF  ( .d(
        \prgm_register/or_signal [360]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[360]) );
  d_ff \prgm_register/genblk1[359].single_DFF  ( .d(
        \prgm_register/or_signal [359]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[359]) );
  d_ff \prgm_register/genblk1[358].single_DFF  ( .d(
        \prgm_register/or_signal [358]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[358]) );
  d_ff \prgm_register/genblk1[357].single_DFF  ( .d(
        \prgm_register/or_signal [357]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[357]) );
  d_ff \prgm_register/genblk1[356].single_DFF  ( .d(
        \prgm_register/or_signal [356]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[356]) );
  d_ff \prgm_register/genblk1[355].single_DFF  ( .d(
        \prgm_register/or_signal [355]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[355]) );
  d_ff \prgm_register/genblk1[354].single_DFF  ( .d(
        \prgm_register/or_signal [354]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[354]) );
  d_ff \prgm_register/genblk1[353].single_DFF  ( .d(
        \prgm_register/or_signal [353]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[353]) );
  d_ff \prgm_register/genblk1[352].single_DFF  ( .d(
        \prgm_register/or_signal [352]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[352]) );
  d_ff \prgm_register/genblk1[351].single_DFF  ( .d(
        \prgm_register/or_signal [351]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[351]) );
  d_ff \prgm_register/genblk1[350].single_DFF  ( .d(
        \prgm_register/or_signal [350]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[350]) );
  d_ff \prgm_register/genblk1[349].single_DFF  ( .d(
        \prgm_register/or_signal [349]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[349]) );
  d_ff \prgm_register/genblk1[348].single_DFF  ( .d(
        \prgm_register/or_signal [348]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[348]) );
  d_ff \prgm_register/genblk1[347].single_DFF  ( .d(
        \prgm_register/or_signal [347]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[347]) );
  d_ff \prgm_register/genblk1[346].single_DFF  ( .d(
        \prgm_register/or_signal [346]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[346]) );
  d_ff \prgm_register/genblk1[345].single_DFF  ( .d(
        \prgm_register/or_signal [345]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[345]) );
  d_ff \prgm_register/genblk1[344].single_DFF  ( .d(
        \prgm_register/or_signal [344]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[344]) );
  d_ff \prgm_register/genblk1[343].single_DFF  ( .d(
        \prgm_register/or_signal [343]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[343]) );
  d_ff \prgm_register/genblk1[342].single_DFF  ( .d(
        \prgm_register/or_signal [342]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[342]) );
  d_ff \prgm_register/genblk1[341].single_DFF  ( .d(
        \prgm_register/or_signal [341]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[341]) );
  d_ff \prgm_register/genblk1[340].single_DFF  ( .d(
        \prgm_register/or_signal [340]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[340]) );
  d_ff \prgm_register/genblk1[339].single_DFF  ( .d(
        \prgm_register/or_signal [339]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[339]) );
  d_ff \prgm_register/genblk1[338].single_DFF  ( .d(
        \prgm_register/or_signal [338]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[338]) );
  d_ff \prgm_register/genblk1[337].single_DFF  ( .d(
        \prgm_register/or_signal [337]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[337]) );
  d_ff \prgm_register/genblk1[336].single_DFF  ( .d(
        \prgm_register/or_signal [336]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[336]) );
  d_ff \prgm_register/genblk1[335].single_DFF  ( .d(
        \prgm_register/or_signal [335]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[335]) );
  d_ff \prgm_register/genblk1[334].single_DFF  ( .d(
        \prgm_register/or_signal [334]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[334]) );
  d_ff \prgm_register/genblk1[333].single_DFF  ( .d(
        \prgm_register/or_signal [333]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[333]) );
  d_ff \prgm_register/genblk1[332].single_DFF  ( .d(
        \prgm_register/or_signal [332]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[332]) );
  d_ff \prgm_register/genblk1[331].single_DFF  ( .d(
        \prgm_register/or_signal [331]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[331]) );
  d_ff \prgm_register/genblk1[330].single_DFF  ( .d(
        \prgm_register/or_signal [330]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[330]) );
  d_ff \prgm_register/genblk1[329].single_DFF  ( .d(
        \prgm_register/or_signal [329]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[329]) );
  d_ff \prgm_register/genblk1[328].single_DFF  ( .d(
        \prgm_register/or_signal [328]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[328]) );
  d_ff \prgm_register/genblk1[327].single_DFF  ( .d(
        \prgm_register/or_signal [327]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[327]) );
  d_ff \prgm_register/genblk1[326].single_DFF  ( .d(
        \prgm_register/or_signal [326]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[326]) );
  d_ff \prgm_register/genblk1[325].single_DFF  ( .d(
        \prgm_register/or_signal [325]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[325]) );
  d_ff \prgm_register/genblk1[324].single_DFF  ( .d(
        \prgm_register/or_signal [324]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[324]) );
  d_ff \prgm_register/genblk1[323].single_DFF  ( .d(
        \prgm_register/or_signal [323]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[323]) );
  d_ff \prgm_register/genblk1[322].single_DFF  ( .d(
        \prgm_register/or_signal [322]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[322]) );
  d_ff \prgm_register/genblk1[321].single_DFF  ( .d(
        \prgm_register/or_signal [321]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[321]) );
  d_ff \prgm_register/genblk1[320].single_DFF  ( .d(
        \prgm_register/or_signal [320]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[320]) );
  d_ff \prgm_register/genblk1[319].single_DFF  ( .d(
        \prgm_register/or_signal [319]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[319]) );
  d_ff \prgm_register/genblk1[318].single_DFF  ( .d(
        \prgm_register/or_signal [318]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[318]) );
  d_ff \prgm_register/genblk1[317].single_DFF  ( .d(
        \prgm_register/or_signal [317]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[317]) );
  d_ff \prgm_register/genblk1[316].single_DFF  ( .d(
        \prgm_register/or_signal [316]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[316]) );
  d_ff \prgm_register/genblk1[315].single_DFF  ( .d(
        \prgm_register/or_signal [315]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[315]) );
  d_ff \prgm_register/genblk1[314].single_DFF  ( .d(
        \prgm_register/or_signal [314]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[314]) );
  d_ff \prgm_register/genblk1[313].single_DFF  ( .d(
        \prgm_register/or_signal [313]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[313]) );
  d_ff \prgm_register/genblk1[312].single_DFF  ( .d(
        \prgm_register/or_signal [312]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[312]) );
  d_ff \prgm_register/genblk1[311].single_DFF  ( .d(
        \prgm_register/or_signal [311]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[311]) );
  d_ff \prgm_register/genblk1[310].single_DFF  ( .d(
        \prgm_register/or_signal [310]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[310]) );
  d_ff \prgm_register/genblk1[309].single_DFF  ( .d(
        \prgm_register/or_signal [309]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[309]) );
  d_ff \prgm_register/genblk1[308].single_DFF  ( .d(
        \prgm_register/or_signal [308]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[308]) );
  d_ff \prgm_register/genblk1[307].single_DFF  ( .d(
        \prgm_register/or_signal [307]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[307]) );
  d_ff \prgm_register/genblk1[306].single_DFF  ( .d(
        \prgm_register/or_signal [306]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[306]) );
  d_ff \prgm_register/genblk1[305].single_DFF  ( .d(
        \prgm_register/or_signal [305]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[305]) );
  d_ff \prgm_register/genblk1[304].single_DFF  ( .d(
        \prgm_register/or_signal [304]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[304]) );
  d_ff \prgm_register/genblk1[303].single_DFF  ( .d(
        \prgm_register/or_signal [303]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[303]) );
  d_ff \prgm_register/genblk1[302].single_DFF  ( .d(
        \prgm_register/or_signal [302]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[302]) );
  d_ff \prgm_register/genblk1[301].single_DFF  ( .d(
        \prgm_register/or_signal [301]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[301]) );
  d_ff \prgm_register/genblk1[300].single_DFF  ( .d(
        \prgm_register/or_signal [300]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[300]) );
  d_ff \prgm_register/genblk1[299].single_DFF  ( .d(
        \prgm_register/or_signal [299]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[299]) );
  d_ff \prgm_register/genblk1[298].single_DFF  ( .d(
        \prgm_register/or_signal [298]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[298]) );
  d_ff \prgm_register/genblk1[297].single_DFF  ( .d(
        \prgm_register/or_signal [297]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[297]) );
  d_ff \prgm_register/genblk1[296].single_DFF  ( .d(
        \prgm_register/or_signal [296]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[296]) );
  d_ff \prgm_register/genblk1[295].single_DFF  ( .d(
        \prgm_register/or_signal [295]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[295]) );
  d_ff \prgm_register/genblk1[294].single_DFF  ( .d(
        \prgm_register/or_signal [294]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[294]) );
  d_ff \prgm_register/genblk1[293].single_DFF  ( .d(
        \prgm_register/or_signal [293]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[293]) );
  d_ff \prgm_register/genblk1[292].single_DFF  ( .d(
        \prgm_register/or_signal [292]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[292]) );
  d_ff \prgm_register/genblk1[291].single_DFF  ( .d(
        \prgm_register/or_signal [291]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[291]) );
  d_ff \prgm_register/genblk1[290].single_DFF  ( .d(
        \prgm_register/or_signal [290]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[290]) );
  d_ff \prgm_register/genblk1[289].single_DFF  ( .d(
        \prgm_register/or_signal [289]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[289]) );
  d_ff \prgm_register/genblk1[288].single_DFF  ( .d(
        \prgm_register/or_signal [288]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[288]) );
  d_ff \prgm_register/genblk1[287].single_DFF  ( .d(
        \prgm_register/or_signal [287]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[287]) );
  d_ff \prgm_register/genblk1[286].single_DFF  ( .d(
        \prgm_register/or_signal [286]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[286]) );
  d_ff \prgm_register/genblk1[285].single_DFF  ( .d(
        \prgm_register/or_signal [285]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[285]) );
  d_ff \prgm_register/genblk1[284].single_DFF  ( .d(
        \prgm_register/or_signal [284]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[284]) );
  d_ff \prgm_register/genblk1[283].single_DFF  ( .d(
        \prgm_register/or_signal [283]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[283]) );
  d_ff \prgm_register/genblk1[282].single_DFF  ( .d(
        \prgm_register/or_signal [282]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[282]) );
  d_ff \prgm_register/genblk1[281].single_DFF  ( .d(
        \prgm_register/or_signal [281]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[281]) );
  d_ff \prgm_register/genblk1[280].single_DFF  ( .d(
        \prgm_register/or_signal [280]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[280]) );
  d_ff \prgm_register/genblk1[279].single_DFF  ( .d(
        \prgm_register/or_signal [279]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[279]) );
  d_ff \prgm_register/genblk1[278].single_DFF  ( .d(
        \prgm_register/or_signal [278]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[278]) );
  d_ff \prgm_register/genblk1[277].single_DFF  ( .d(
        \prgm_register/or_signal [277]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[277]) );
  d_ff \prgm_register/genblk1[276].single_DFF  ( .d(
        \prgm_register/or_signal [276]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[276]) );
  d_ff \prgm_register/genblk1[275].single_DFF  ( .d(
        \prgm_register/or_signal [275]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[275]) );
  d_ff \prgm_register/genblk1[274].single_DFF  ( .d(
        \prgm_register/or_signal [274]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[274]) );
  d_ff \prgm_register/genblk1[273].single_DFF  ( .d(
        \prgm_register/or_signal [273]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[273]) );
  d_ff \prgm_register/genblk1[272].single_DFF  ( .d(
        \prgm_register/or_signal [272]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[272]) );
  d_ff \prgm_register/genblk1[271].single_DFF  ( .d(
        \prgm_register/or_signal [271]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[271]) );
  d_ff \prgm_register/genblk1[270].single_DFF  ( .d(
        \prgm_register/or_signal [270]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[270]) );
  d_ff \prgm_register/genblk1[269].single_DFF  ( .d(
        \prgm_register/or_signal [269]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[269]) );
  d_ff \prgm_register/genblk1[268].single_DFF  ( .d(
        \prgm_register/or_signal [268]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[268]) );
  d_ff \prgm_register/genblk1[267].single_DFF  ( .d(
        \prgm_register/or_signal [267]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[267]) );
  d_ff \prgm_register/genblk1[266].single_DFF  ( .d(
        \prgm_register/or_signal [266]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[266]) );
  d_ff \prgm_register/genblk1[265].single_DFF  ( .d(
        \prgm_register/or_signal [265]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[265]) );
  d_ff \prgm_register/genblk1[264].single_DFF  ( .d(
        \prgm_register/or_signal [264]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[264]) );
  d_ff \prgm_register/genblk1[263].single_DFF  ( .d(
        \prgm_register/or_signal [263]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[263]) );
  d_ff \prgm_register/genblk1[262].single_DFF  ( .d(
        \prgm_register/or_signal [262]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[262]) );
  d_ff \prgm_register/genblk1[261].single_DFF  ( .d(
        \prgm_register/or_signal [261]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[261]) );
  d_ff \prgm_register/genblk1[260].single_DFF  ( .d(
        \prgm_register/or_signal [260]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[260]) );
  d_ff \prgm_register/genblk1[259].single_DFF  ( .d(
        \prgm_register/or_signal [259]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[259]) );
  d_ff \prgm_register/genblk1[258].single_DFF  ( .d(
        \prgm_register/or_signal [258]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[258]) );
  d_ff \prgm_register/genblk1[257].single_DFF  ( .d(
        \prgm_register/or_signal [257]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[257]) );
  d_ff \prgm_register/genblk1[256].single_DFF  ( .d(
        \prgm_register/or_signal [256]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[256]) );
  d_ff \prgm_register/genblk1[255].single_DFF  ( .d(
        \prgm_register/or_signal [255]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[255]) );
  d_ff \prgm_register/genblk1[254].single_DFF  ( .d(
        \prgm_register/or_signal [254]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[254]) );
  d_ff \prgm_register/genblk1[253].single_DFF  ( .d(
        \prgm_register/or_signal [253]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[253]) );
  d_ff \prgm_register/genblk1[252].single_DFF  ( .d(
        \prgm_register/or_signal [252]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[252]) );
  d_ff \prgm_register/genblk1[251].single_DFF  ( .d(
        \prgm_register/or_signal [251]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[251]) );
  d_ff \prgm_register/genblk1[250].single_DFF  ( .d(
        \prgm_register/or_signal [250]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[250]) );
  d_ff \prgm_register/genblk1[249].single_DFF  ( .d(
        \prgm_register/or_signal [249]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[249]) );
  d_ff \prgm_register/genblk1[248].single_DFF  ( .d(
        \prgm_register/or_signal [248]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[248]) );
  d_ff \prgm_register/genblk1[247].single_DFF  ( .d(
        \prgm_register/or_signal [247]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[247]) );
  d_ff \prgm_register/genblk1[246].single_DFF  ( .d(
        \prgm_register/or_signal [246]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[246]) );
  d_ff \prgm_register/genblk1[245].single_DFF  ( .d(
        \prgm_register/or_signal [245]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[245]) );
  d_ff \prgm_register/genblk1[244].single_DFF  ( .d(
        \prgm_register/or_signal [244]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[244]) );
  d_ff \prgm_register/genblk1[243].single_DFF  ( .d(
        \prgm_register/or_signal [243]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[243]) );
  d_ff \prgm_register/genblk1[242].single_DFF  ( .d(
        \prgm_register/or_signal [242]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[242]) );
  d_ff \prgm_register/genblk1[241].single_DFF  ( .d(
        \prgm_register/or_signal [241]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[241]) );
  d_ff \prgm_register/genblk1[240].single_DFF  ( .d(
        \prgm_register/or_signal [240]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[240]) );
  d_ff \prgm_register/genblk1[239].single_DFF  ( .d(
        \prgm_register/or_signal [239]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[239]) );
  d_ff \prgm_register/genblk1[238].single_DFF  ( .d(
        \prgm_register/or_signal [238]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[238]) );
  d_ff \prgm_register/genblk1[237].single_DFF  ( .d(
        \prgm_register/or_signal [237]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[237]) );
  d_ff \prgm_register/genblk1[236].single_DFF  ( .d(
        \prgm_register/or_signal [236]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[236]) );
  d_ff \prgm_register/genblk1[235].single_DFF  ( .d(
        \prgm_register/or_signal [235]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[235]) );
  d_ff \prgm_register/genblk1[234].single_DFF  ( .d(
        \prgm_register/or_signal [234]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[234]) );
  d_ff \prgm_register/genblk1[233].single_DFF  ( .d(
        \prgm_register/or_signal [233]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[233]) );
  d_ff \prgm_register/genblk1[232].single_DFF  ( .d(
        \prgm_register/or_signal [232]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[232]) );
  d_ff \prgm_register/genblk1[231].single_DFF  ( .d(
        \prgm_register/or_signal [231]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[231]) );
  d_ff \prgm_register/genblk1[230].single_DFF  ( .d(
        \prgm_register/or_signal [230]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[230]) );
  d_ff \prgm_register/genblk1[229].single_DFF  ( .d(
        \prgm_register/or_signal [229]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[229]) );
  d_ff \prgm_register/genblk1[228].single_DFF  ( .d(
        \prgm_register/or_signal [228]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[228]) );
  d_ff \prgm_register/genblk1[227].single_DFF  ( .d(
        \prgm_register/or_signal [227]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[227]) );
  d_ff \prgm_register/genblk1[226].single_DFF  ( .d(
        \prgm_register/or_signal [226]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[226]) );
  d_ff \prgm_register/genblk1[225].single_DFF  ( .d(
        \prgm_register/or_signal [225]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[225]) );
  d_ff \prgm_register/genblk1[224].single_DFF  ( .d(
        \prgm_register/or_signal [224]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[224]) );
  d_ff \prgm_register/genblk1[223].single_DFF  ( .d(
        \prgm_register/or_signal [223]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[223]) );
  d_ff \prgm_register/genblk1[222].single_DFF  ( .d(
        \prgm_register/or_signal [222]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[222]) );
  d_ff \prgm_register/genblk1[221].single_DFF  ( .d(
        \prgm_register/or_signal [221]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[221]) );
  d_ff \prgm_register/genblk1[220].single_DFF  ( .d(
        \prgm_register/or_signal [220]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[220]) );
  d_ff \prgm_register/genblk1[219].single_DFF  ( .d(
        \prgm_register/or_signal [219]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[219]) );
  d_ff \prgm_register/genblk1[218].single_DFF  ( .d(
        \prgm_register/or_signal [218]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[218]) );
  d_ff \prgm_register/genblk1[217].single_DFF  ( .d(
        \prgm_register/or_signal [217]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[217]) );
  d_ff \prgm_register/genblk1[216].single_DFF  ( .d(
        \prgm_register/or_signal [216]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[216]) );
  d_ff \prgm_register/genblk1[215].single_DFF  ( .d(
        \prgm_register/or_signal [215]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[215]) );
  d_ff \prgm_register/genblk1[214].single_DFF  ( .d(
        \prgm_register/or_signal [214]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[214]) );
  d_ff \prgm_register/genblk1[213].single_DFF  ( .d(
        \prgm_register/or_signal [213]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[213]) );
  d_ff \prgm_register/genblk1[212].single_DFF  ( .d(
        \prgm_register/or_signal [212]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[212]) );
  d_ff \prgm_register/genblk1[211].single_DFF  ( .d(
        \prgm_register/or_signal [211]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[211]) );
  d_ff \prgm_register/genblk1[210].single_DFF  ( .d(
        \prgm_register/or_signal [210]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[210]) );
  d_ff \prgm_register/genblk1[209].single_DFF  ( .d(
        \prgm_register/or_signal [209]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[209]) );
  d_ff \prgm_register/genblk1[208].single_DFF  ( .d(
        \prgm_register/or_signal [208]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[208]) );
  d_ff \prgm_register/genblk1[207].single_DFF  ( .d(
        \prgm_register/or_signal [207]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[207]) );
  d_ff \prgm_register/genblk1[206].single_DFF  ( .d(
        \prgm_register/or_signal [206]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[206]) );
  d_ff \prgm_register/genblk1[205].single_DFF  ( .d(
        \prgm_register/or_signal [205]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[205]) );
  d_ff \prgm_register/genblk1[204].single_DFF  ( .d(
        \prgm_register/or_signal [204]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[204]) );
  d_ff \prgm_register/genblk1[203].single_DFF  ( .d(
        \prgm_register/or_signal [203]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[203]) );
  d_ff \prgm_register/genblk1[202].single_DFF  ( .d(
        \prgm_register/or_signal [202]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[202]) );
  d_ff \prgm_register/genblk1[201].single_DFF  ( .d(
        \prgm_register/or_signal [201]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[201]) );
  d_ff \prgm_register/genblk1[200].single_DFF  ( .d(
        \prgm_register/or_signal [200]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[200]) );
  d_ff \prgm_register/genblk1[199].single_DFF  ( .d(
        \prgm_register/or_signal [199]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[199]) );
  d_ff \prgm_register/genblk1[198].single_DFF  ( .d(
        \prgm_register/or_signal [198]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[198]) );
  d_ff \prgm_register/genblk1[197].single_DFF  ( .d(
        \prgm_register/or_signal [197]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[197]) );
  d_ff \prgm_register/genblk1[196].single_DFF  ( .d(
        \prgm_register/or_signal [196]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[196]) );
  d_ff \prgm_register/genblk1[195].single_DFF  ( .d(
        \prgm_register/or_signal [195]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[195]) );
  d_ff \prgm_register/genblk1[194].single_DFF  ( .d(
        \prgm_register/or_signal [194]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[194]) );
  d_ff \prgm_register/genblk1[193].single_DFF  ( .d(
        \prgm_register/or_signal [193]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[193]) );
  d_ff \prgm_register/genblk1[192].single_DFF  ( .d(
        \prgm_register/or_signal [192]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[192]) );
  d_ff \prgm_register/genblk1[191].single_DFF  ( .d(
        \prgm_register/or_signal [191]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[191]) );
  d_ff \prgm_register/genblk1[190].single_DFF  ( .d(
        \prgm_register/or_signal [190]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[190]) );
  d_ff \prgm_register/genblk1[189].single_DFF  ( .d(
        \prgm_register/or_signal [189]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[189]) );
  d_ff \prgm_register/genblk1[188].single_DFF  ( .d(
        \prgm_register/or_signal [188]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[188]) );
  d_ff \prgm_register/genblk1[187].single_DFF  ( .d(
        \prgm_register/or_signal [187]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[187]) );
  d_ff \prgm_register/genblk1[186].single_DFF  ( .d(
        \prgm_register/or_signal [186]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[186]) );
  d_ff \prgm_register/genblk1[185].single_DFF  ( .d(
        \prgm_register/or_signal [185]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[185]) );
  d_ff \prgm_register/genblk1[184].single_DFF  ( .d(
        \prgm_register/or_signal [184]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[184]) );
  d_ff \prgm_register/genblk1[183].single_DFF  ( .d(
        \prgm_register/or_signal [183]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[183]) );
  d_ff \prgm_register/genblk1[182].single_DFF  ( .d(
        \prgm_register/or_signal [182]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[182]) );
  d_ff \prgm_register/genblk1[181].single_DFF  ( .d(
        \prgm_register/or_signal [181]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[181]) );
  d_ff \prgm_register/genblk1[180].single_DFF  ( .d(
        \prgm_register/or_signal [180]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[180]) );
  d_ff \prgm_register/genblk1[179].single_DFF  ( .d(
        \prgm_register/or_signal [179]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[179]) );
  d_ff \prgm_register/genblk1[178].single_DFF  ( .d(
        \prgm_register/or_signal [178]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[178]) );
  d_ff \prgm_register/genblk1[177].single_DFF  ( .d(
        \prgm_register/or_signal [177]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[177]) );
  d_ff \prgm_register/genblk1[176].single_DFF  ( .d(
        \prgm_register/or_signal [176]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[176]) );
  d_ff \prgm_register/genblk1[175].single_DFF  ( .d(
        \prgm_register/or_signal [175]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[175]) );
  d_ff \prgm_register/genblk1[174].single_DFF  ( .d(
        \prgm_register/or_signal [174]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[174]) );
  d_ff \prgm_register/genblk1[173].single_DFF  ( .d(
        \prgm_register/or_signal [173]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[173]) );
  d_ff \prgm_register/genblk1[172].single_DFF  ( .d(
        \prgm_register/or_signal [172]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[172]) );
  d_ff \prgm_register/genblk1[171].single_DFF  ( .d(
        \prgm_register/or_signal [171]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[171]) );
  d_ff \prgm_register/genblk1[170].single_DFF  ( .d(
        \prgm_register/or_signal [170]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[170]) );
  d_ff \prgm_register/genblk1[169].single_DFF  ( .d(
        \prgm_register/or_signal [169]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[169]) );
  d_ff \prgm_register/genblk1[168].single_DFF  ( .d(
        \prgm_register/or_signal [168]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[168]) );
  d_ff \prgm_register/genblk1[167].single_DFF  ( .d(
        \prgm_register/or_signal [167]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[167]) );
  d_ff \prgm_register/genblk1[166].single_DFF  ( .d(
        \prgm_register/or_signal [166]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[166]) );
  d_ff \prgm_register/genblk1[165].single_DFF  ( .d(
        \prgm_register/or_signal [165]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[165]) );
  d_ff \prgm_register/genblk1[164].single_DFF  ( .d(
        \prgm_register/or_signal [164]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[164]) );
  d_ff \prgm_register/genblk1[163].single_DFF  ( .d(
        \prgm_register/or_signal [163]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[163]) );
  d_ff \prgm_register/genblk1[162].single_DFF  ( .d(
        \prgm_register/or_signal [162]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[162]) );
  d_ff \prgm_register/genblk1[161].single_DFF  ( .d(
        \prgm_register/or_signal [161]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[161]) );
  d_ff \prgm_register/genblk1[160].single_DFF  ( .d(
        \prgm_register/or_signal [160]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[160]) );
  d_ff \prgm_register/genblk1[159].single_DFF  ( .d(
        \prgm_register/or_signal [159]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[159]) );
  d_ff \prgm_register/genblk1[158].single_DFF  ( .d(
        \prgm_register/or_signal [158]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[158]) );
  d_ff \prgm_register/genblk1[157].single_DFF  ( .d(
        \prgm_register/or_signal [157]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[157]) );
  d_ff \prgm_register/genblk1[156].single_DFF  ( .d(
        \prgm_register/or_signal [156]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[156]) );
  d_ff \prgm_register/genblk1[155].single_DFF  ( .d(
        \prgm_register/or_signal [155]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[155]) );
  d_ff \prgm_register/genblk1[154].single_DFF  ( .d(
        \prgm_register/or_signal [154]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[154]) );
  d_ff \prgm_register/genblk1[153].single_DFF  ( .d(
        \prgm_register/or_signal [153]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[153]) );
  d_ff \prgm_register/genblk1[152].single_DFF  ( .d(
        \prgm_register/or_signal [152]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[152]) );
  d_ff \prgm_register/genblk1[151].single_DFF  ( .d(
        \prgm_register/or_signal [151]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[151]) );
  d_ff \prgm_register/genblk1[150].single_DFF  ( .d(
        \prgm_register/or_signal [150]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[150]) );
  d_ff \prgm_register/genblk1[149].single_DFF  ( .d(
        \prgm_register/or_signal [149]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[149]) );
  d_ff \prgm_register/genblk1[148].single_DFF  ( .d(
        \prgm_register/or_signal [148]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[148]) );
  d_ff \prgm_register/genblk1[147].single_DFF  ( .d(
        \prgm_register/or_signal [147]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[147]) );
  d_ff \prgm_register/genblk1[146].single_DFF  ( .d(
        \prgm_register/or_signal [146]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[146]) );
  d_ff \prgm_register/genblk1[145].single_DFF  ( .d(
        \prgm_register/or_signal [145]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[145]) );
  d_ff \prgm_register/genblk1[144].single_DFF  ( .d(
        \prgm_register/or_signal [144]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[144]) );
  d_ff \prgm_register/genblk1[143].single_DFF  ( .d(
        \prgm_register/or_signal [143]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[143]) );
  d_ff \prgm_register/genblk1[142].single_DFF  ( .d(
        \prgm_register/or_signal [142]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[142]) );
  d_ff \prgm_register/genblk1[141].single_DFF  ( .d(
        \prgm_register/or_signal [141]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[141]) );
  d_ff \prgm_register/genblk1[140].single_DFF  ( .d(
        \prgm_register/or_signal [140]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[140]) );
  d_ff \prgm_register/genblk1[139].single_DFF  ( .d(
        \prgm_register/or_signal [139]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[139]) );
  d_ff \prgm_register/genblk1[138].single_DFF  ( .d(
        \prgm_register/or_signal [138]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[138]) );
  d_ff \prgm_register/genblk1[137].single_DFF  ( .d(
        \prgm_register/or_signal [137]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[137]) );
  d_ff \prgm_register/genblk1[136].single_DFF  ( .d(
        \prgm_register/or_signal [136]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[136]) );
  d_ff \prgm_register/genblk1[135].single_DFF  ( .d(
        \prgm_register/or_signal [135]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[135]) );
  d_ff \prgm_register/genblk1[134].single_DFF  ( .d(
        \prgm_register/or_signal [134]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[134]) );
  d_ff \prgm_register/genblk1[133].single_DFF  ( .d(
        \prgm_register/or_signal [133]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[133]) );
  d_ff \prgm_register/genblk1[132].single_DFF  ( .d(
        \prgm_register/or_signal [132]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[132]) );
  d_ff \prgm_register/genblk1[131].single_DFF  ( .d(
        \prgm_register/or_signal [131]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[131]) );
  d_ff \prgm_register/genblk1[130].single_DFF  ( .d(
        \prgm_register/or_signal [130]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[130]) );
  d_ff \prgm_register/genblk1[129].single_DFF  ( .d(
        \prgm_register/or_signal [129]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[129]) );
  d_ff \prgm_register/genblk1[128].single_DFF  ( .d(
        \prgm_register/or_signal [128]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[128]) );
  d_ff \prgm_register/genblk1[127].single_DFF  ( .d(
        \prgm_register/or_signal [127]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[127]) );
  d_ff \prgm_register/genblk1[126].single_DFF  ( .d(
        \prgm_register/or_signal [126]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[126]) );
  d_ff \prgm_register/genblk1[125].single_DFF  ( .d(
        \prgm_register/or_signal [125]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[125]) );
  d_ff \prgm_register/genblk1[124].single_DFF  ( .d(
        \prgm_register/or_signal [124]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[124]) );
  d_ff \prgm_register/genblk1[123].single_DFF  ( .d(
        \prgm_register/or_signal [123]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[123]) );
  d_ff \prgm_register/genblk1[122].single_DFF  ( .d(
        \prgm_register/or_signal [122]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[122]) );
  d_ff \prgm_register/genblk1[121].single_DFF  ( .d(
        \prgm_register/or_signal [121]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[121]) );
  d_ff \prgm_register/genblk1[120].single_DFF  ( .d(
        \prgm_register/or_signal [120]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[120]) );
  d_ff \prgm_register/genblk1[119].single_DFF  ( .d(
        \prgm_register/or_signal [119]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[119]) );
  d_ff \prgm_register/genblk1[118].single_DFF  ( .d(
        \prgm_register/or_signal [118]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[118]) );
  d_ff \prgm_register/genblk1[117].single_DFF  ( .d(
        \prgm_register/or_signal [117]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[117]) );
  d_ff \prgm_register/genblk1[116].single_DFF  ( .d(
        \prgm_register/or_signal [116]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[116]) );
  d_ff \prgm_register/genblk1[115].single_DFF  ( .d(
        \prgm_register/or_signal [115]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[115]) );
  d_ff \prgm_register/genblk1[114].single_DFF  ( .d(
        \prgm_register/or_signal [114]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[114]) );
  d_ff \prgm_register/genblk1[113].single_DFF  ( .d(
        \prgm_register/or_signal [113]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[113]) );
  d_ff \prgm_register/genblk1[112].single_DFF  ( .d(
        \prgm_register/or_signal [112]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[112]) );
  d_ff \prgm_register/genblk1[111].single_DFF  ( .d(
        \prgm_register/or_signal [111]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[111]) );
  d_ff \prgm_register/genblk1[110].single_DFF  ( .d(
        \prgm_register/or_signal [110]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[110]) );
  d_ff \prgm_register/genblk1[109].single_DFF  ( .d(
        \prgm_register/or_signal [109]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[109]) );
  d_ff \prgm_register/genblk1[108].single_DFF  ( .d(
        \prgm_register/or_signal [108]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[108]) );
  d_ff \prgm_register/genblk1[107].single_DFF  ( .d(
        \prgm_register/or_signal [107]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[107]) );
  d_ff \prgm_register/genblk1[106].single_DFF  ( .d(
        \prgm_register/or_signal [106]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[106]) );
  d_ff \prgm_register/genblk1[105].single_DFF  ( .d(
        \prgm_register/or_signal [105]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[105]) );
  d_ff \prgm_register/genblk1[104].single_DFF  ( .d(
        \prgm_register/or_signal [104]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[104]) );
  d_ff \prgm_register/genblk1[103].single_DFF  ( .d(
        \prgm_register/or_signal [103]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[103]) );
  d_ff \prgm_register/genblk1[102].single_DFF  ( .d(
        \prgm_register/or_signal [102]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[102]) );
  d_ff \prgm_register/genblk1[101].single_DFF  ( .d(
        \prgm_register/or_signal [101]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[101]) );
  d_ff \prgm_register/genblk1[100].single_DFF  ( .d(
        \prgm_register/or_signal [100]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[100]) );
  d_ff \prgm_register/genblk1[99].single_DFF  ( .d(
        \prgm_register/or_signal [99]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[99]) );
  d_ff \prgm_register/genblk1[98].single_DFF  ( .d(
        \prgm_register/or_signal [98]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[98]) );
  d_ff \prgm_register/genblk1[97].single_DFF  ( .d(
        \prgm_register/or_signal [97]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[97]) );
  d_ff \prgm_register/genblk1[96].single_DFF  ( .d(
        \prgm_register/or_signal [96]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[96]) );
  d_ff \prgm_register/genblk1[95].single_DFF  ( .d(
        \prgm_register/or_signal [95]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[95]) );
  d_ff \prgm_register/genblk1[94].single_DFF  ( .d(
        \prgm_register/or_signal [94]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[94]) );
  d_ff \prgm_register/genblk1[93].single_DFF  ( .d(
        \prgm_register/or_signal [93]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[93]) );
  d_ff \prgm_register/genblk1[92].single_DFF  ( .d(
        \prgm_register/or_signal [92]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[92]) );
  d_ff \prgm_register/genblk1[91].single_DFF  ( .d(
        \prgm_register/or_signal [91]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[91]) );
  d_ff \prgm_register/genblk1[90].single_DFF  ( .d(
        \prgm_register/or_signal [90]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[90]) );
  d_ff \prgm_register/genblk1[89].single_DFF  ( .d(
        \prgm_register/or_signal [89]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[89]) );
  d_ff \prgm_register/genblk1[88].single_DFF  ( .d(
        \prgm_register/or_signal [88]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[88]) );
  d_ff \prgm_register/genblk1[87].single_DFF  ( .d(
        \prgm_register/or_signal [87]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[87]) );
  d_ff \prgm_register/genblk1[86].single_DFF  ( .d(
        \prgm_register/or_signal [86]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[86]) );
  d_ff \prgm_register/genblk1[85].single_DFF  ( .d(
        \prgm_register/or_signal [85]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[85]) );
  d_ff \prgm_register/genblk1[84].single_DFF  ( .d(
        \prgm_register/or_signal [84]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[84]) );
  d_ff \prgm_register/genblk1[83].single_DFF  ( .d(
        \prgm_register/or_signal [83]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[83]) );
  d_ff \prgm_register/genblk1[82].single_DFF  ( .d(
        \prgm_register/or_signal [82]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[82]) );
  d_ff \prgm_register/genblk1[81].single_DFF  ( .d(
        \prgm_register/or_signal [81]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[81]) );
  d_ff \prgm_register/genblk1[80].single_DFF  ( .d(
        \prgm_register/or_signal [80]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[80]) );
  d_ff \prgm_register/genblk1[79].single_DFF  ( .d(
        \prgm_register/or_signal [79]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[79]) );
  d_ff \prgm_register/genblk1[78].single_DFF  ( .d(
        \prgm_register/or_signal [78]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[78]) );
  d_ff \prgm_register/genblk1[77].single_DFF  ( .d(
        \prgm_register/or_signal [77]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[77]) );
  d_ff \prgm_register/genblk1[76].single_DFF  ( .d(
        \prgm_register/or_signal [76]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[76]) );
  d_ff \prgm_register/genblk1[75].single_DFF  ( .d(
        \prgm_register/or_signal [75]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[75]) );
  d_ff \prgm_register/genblk1[74].single_DFF  ( .d(
        \prgm_register/or_signal [74]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[74]) );
  d_ff \prgm_register/genblk1[73].single_DFF  ( .d(
        \prgm_register/or_signal [73]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[73]) );
  d_ff \prgm_register/genblk1[72].single_DFF  ( .d(
        \prgm_register/or_signal [72]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[72]) );
  d_ff \prgm_register/genblk1[71].single_DFF  ( .d(
        \prgm_register/or_signal [71]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[71]) );
  d_ff \prgm_register/genblk1[70].single_DFF  ( .d(
        \prgm_register/or_signal [70]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[70]) );
  d_ff \prgm_register/genblk1[69].single_DFF  ( .d(
        \prgm_register/or_signal [69]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[69]) );
  d_ff \prgm_register/genblk1[68].single_DFF  ( .d(
        \prgm_register/or_signal [68]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[68]) );
  d_ff \prgm_register/genblk1[67].single_DFF  ( .d(
        \prgm_register/or_signal [67]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[67]) );
  d_ff \prgm_register/genblk1[66].single_DFF  ( .d(
        \prgm_register/or_signal [66]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[66]) );
  d_ff \prgm_register/genblk1[65].single_DFF  ( .d(
        \prgm_register/or_signal [65]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[65]) );
  d_ff \prgm_register/genblk1[64].single_DFF  ( .d(
        \prgm_register/or_signal [64]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[64]) );
  d_ff \prgm_register/genblk1[63].single_DFF  ( .d(
        \prgm_register/or_signal [63]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[63]) );
  d_ff \prgm_register/genblk1[62].single_DFF  ( .d(
        \prgm_register/or_signal [62]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[62]) );
  d_ff \prgm_register/genblk1[61].single_DFF  ( .d(
        \prgm_register/or_signal [61]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[61]) );
  d_ff \prgm_register/genblk1[60].single_DFF  ( .d(
        \prgm_register/or_signal [60]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[60]) );
  d_ff \prgm_register/genblk1[59].single_DFF  ( .d(
        \prgm_register/or_signal [59]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[59]) );
  d_ff \prgm_register/genblk1[58].single_DFF  ( .d(
        \prgm_register/or_signal [58]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[58]) );
  d_ff \prgm_register/genblk1[57].single_DFF  ( .d(
        \prgm_register/or_signal [57]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[57]) );
  d_ff \prgm_register/genblk1[56].single_DFF  ( .d(
        \prgm_register/or_signal [56]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[56]) );
  d_ff \prgm_register/genblk1[55].single_DFF  ( .d(
        \prgm_register/or_signal [55]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[55]) );
  d_ff \prgm_register/genblk1[54].single_DFF  ( .d(
        \prgm_register/or_signal [54]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[54]) );
  d_ff \prgm_register/genblk1[53].single_DFF  ( .d(
        \prgm_register/or_signal [53]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[53]) );
  d_ff \prgm_register/genblk1[52].single_DFF  ( .d(
        \prgm_register/or_signal [52]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[52]) );
  d_ff \prgm_register/genblk1[51].single_DFF  ( .d(
        \prgm_register/or_signal [51]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[51]) );
  d_ff \prgm_register/genblk1[50].single_DFF  ( .d(
        \prgm_register/or_signal [50]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[50]) );
  d_ff \prgm_register/genblk1[49].single_DFF  ( .d(
        \prgm_register/or_signal [49]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[49]) );
  d_ff \prgm_register/genblk1[48].single_DFF  ( .d(
        \prgm_register/or_signal [48]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[48]) );
  d_ff \prgm_register/genblk1[47].single_DFF  ( .d(
        \prgm_register/or_signal [47]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[47]) );
  d_ff \prgm_register/genblk1[46].single_DFF  ( .d(
        \prgm_register/or_signal [46]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[46]) );
  d_ff \prgm_register/genblk1[45].single_DFF  ( .d(
        \prgm_register/or_signal [45]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[45]) );
  d_ff \prgm_register/genblk1[44].single_DFF  ( .d(
        \prgm_register/or_signal [44]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[44]) );
  d_ff \prgm_register/genblk1[43].single_DFF  ( .d(
        \prgm_register/or_signal [43]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[43]) );
  d_ff \prgm_register/genblk1[42].single_DFF  ( .d(
        \prgm_register/or_signal [42]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[42]) );
  d_ff \prgm_register/genblk1[41].single_DFF  ( .d(
        \prgm_register/or_signal [41]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[41]) );
  d_ff \prgm_register/genblk1[40].single_DFF  ( .d(
        \prgm_register/or_signal [40]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[40]) );
  d_ff \prgm_register/genblk1[39].single_DFF  ( .d(
        \prgm_register/or_signal [39]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[39]) );
  d_ff \prgm_register/genblk1[38].single_DFF  ( .d(
        \prgm_register/or_signal [38]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[38]) );
  d_ff \prgm_register/genblk1[37].single_DFF  ( .d(
        \prgm_register/or_signal [37]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[37]) );
  d_ff \prgm_register/genblk1[36].single_DFF  ( .d(
        \prgm_register/or_signal [36]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[36]) );
  d_ff \prgm_register/genblk1[35].single_DFF  ( .d(
        \prgm_register/or_signal [35]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[35]) );
  d_ff \prgm_register/genblk1[34].single_DFF  ( .d(
        \prgm_register/or_signal [34]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[34]) );
  d_ff \prgm_register/genblk1[33].single_DFF  ( .d(
        \prgm_register/or_signal [33]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[33]) );
  d_ff \prgm_register/genblk1[32].single_DFF  ( .d(
        \prgm_register/or_signal [32]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[32]) );
  d_ff \prgm_register/genblk1[31].single_DFF  ( .d(
        \prgm_register/or_signal [31]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[31]) );
  d_ff \prgm_register/genblk1[30].single_DFF  ( .d(
        \prgm_register/or_signal [30]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[30]) );
  d_ff \prgm_register/genblk1[29].single_DFF  ( .d(
        \prgm_register/or_signal [29]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[29]) );
  d_ff \prgm_register/genblk1[28].single_DFF  ( .d(
        \prgm_register/or_signal [28]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[28]) );
  d_ff \prgm_register/genblk1[27].single_DFF  ( .d(
        \prgm_register/or_signal [27]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[27]) );
  d_ff \prgm_register/genblk1[26].single_DFF  ( .d(
        \prgm_register/or_signal [26]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[26]) );
  d_ff \prgm_register/genblk1[25].single_DFF  ( .d(
        \prgm_register/or_signal [25]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[25]) );
  d_ff \prgm_register/genblk1[24].single_DFF  ( .d(
        \prgm_register/or_signal [24]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[24]) );
  d_ff \prgm_register/genblk1[23].single_DFF  ( .d(
        \prgm_register/or_signal [23]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[23]) );
  d_ff \prgm_register/genblk1[22].single_DFF  ( .d(
        \prgm_register/or_signal [22]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[22]) );
  d_ff \prgm_register/genblk1[21].single_DFF  ( .d(
        \prgm_register/or_signal [21]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[21]) );
  d_ff \prgm_register/genblk1[20].single_DFF  ( .d(
        \prgm_register/or_signal [20]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[20]) );
  d_ff \prgm_register/genblk1[19].single_DFF  ( .d(
        \prgm_register/or_signal [19]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[19]) );
  d_ff \prgm_register/genblk1[18].single_DFF  ( .d(
        \prgm_register/or_signal [18]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[18]) );
  d_ff \prgm_register/genblk1[17].single_DFF  ( .d(
        \prgm_register/or_signal [17]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[17]) );
  d_ff \prgm_register/genblk1[16].single_DFF  ( .d(
        \prgm_register/or_signal [16]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[16]) );
  d_ff \prgm_register/genblk1[15].single_DFF  ( .d(
        \prgm_register/or_signal [15]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[15]) );
  d_ff \prgm_register/genblk1[14].single_DFF  ( .d(
        \prgm_register/or_signal [14]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[14]) );
  d_ff \prgm_register/genblk1[13].single_DFF  ( .d(
        \prgm_register/or_signal [13]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[13]) );
  d_ff \prgm_register/genblk1[12].single_DFF  ( .d(
        \prgm_register/or_signal [12]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[12]) );
  d_ff \prgm_register/genblk1[11].single_DFF  ( .d(
        \prgm_register/or_signal [11]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[11]) );
  d_ff \prgm_register/genblk1[10].single_DFF  ( .d(
        \prgm_register/or_signal [10]), .clk(clk), .R(
        \prgm_register/clear_not ), .Q(a[10]) );
  d_ff \prgm_register/genblk1[9].single_DFF  ( .d(\prgm_register/or_signal [9]), 
        .clk(clk), .R(\prgm_register/clear_not ), .Q(a[9]) );
  d_ff \prgm_register/genblk1[8].single_DFF  ( .d(\prgm_register/or_signal [8]), 
        .clk(clk), .R(\prgm_register/clear_not ), .Q(a[8]) );
  d_ff \prgm_register/genblk1[7].single_DFF  ( .d(\prgm_register/or_signal [7]), 
        .clk(clk), .R(\prgm_register/clear_not ), .Q(a[7]) );
  d_ff \prgm_register/genblk1[6].single_DFF  ( .d(\prgm_register/or_signal [6]), 
        .clk(clk), .R(\prgm_register/clear_not ), .Q(a[6]) );
  d_ff \prgm_register/genblk1[5].single_DFF  ( .d(\prgm_register/or_signal [5]), 
        .clk(clk), .R(\prgm_register/clear_not ), .Q(a[5]) );
  d_ff \prgm_register/genblk1[4].single_DFF  ( .d(\prgm_register/or_signal [4]), 
        .clk(clk), .R(\prgm_register/clear_not ), .Q(a[4]) );
  d_ff \prgm_register/genblk1[3].single_DFF  ( .d(\prgm_register/or_signal [3]), 
        .clk(clk), .R(\prgm_register/clear_not ), .Q(a[3]) );
  d_ff \prgm_register/genblk1[2].single_DFF  ( .d(\prgm_register/or_signal [2]), 
        .clk(clk), .R(\prgm_register/clear_not ), .Q(a[2]) );
  d_ff \prgm_register/genblk1[1].single_DFF  ( .d(\prgm_register/or_signal [1]), 
        .clk(clk), .R(\prgm_register/clear_not ), .Q(a[1]) );
  d_ff \prgm_register/first_DFF  ( .d(\prgm_register/or_signal [0]), .clk(clk), 
        .R(\prgm_register/clear_not ), .Q(a[0]) );
  inv \comparator/U2046  ( .a(\comparator/N1 ), .out(\comparator/n2046 ) );
  inv \comparator/U2045  ( .a(\comparator/N0 ), .out(\comparator/n2045 ) );
  inv \comparator/U2044  ( .a(\comparator/N3 ), .out(\comparator/n2044 ) );
  inv \comparator/U2043  ( .a(\comparator/N2 ), .out(\comparator/n2043 ) );
  inv \comparator/U2042  ( .a(\comparator/N5 ), .out(\comparator/n2042 ) );
  inv \comparator/U2041  ( .a(\comparator/N4 ), .out(\comparator/n2041 ) );
  inv \comparator/U2040  ( .a(\comparator/N7 ), .out(\comparator/n2040 ) );
  inv \comparator/U2039  ( .a(\comparator/N6 ), .out(\comparator/n2039 ) );
  inv \comparator/U2038  ( .a(\comparator/N9 ), .out(\comparator/n2038 ) );
  inv \comparator/U2037  ( .a(\comparator/N8 ), .out(\comparator/n2037 ) );
  inv \comparator/U2036  ( .a(\comparator/N11 ), .out(\comparator/n2036 ) );
  inv \comparator/U2035  ( .a(\comparator/N10 ), .out(\comparator/n2035 ) );
  inv \comparator/U2034  ( .a(\comparator/N13 ), .out(\comparator/n2034 ) );
  inv \comparator/U2033  ( .a(\comparator/N12 ), .out(\comparator/n2033 ) );
  inv \comparator/U2032  ( .a(\comparator/N15 ), .out(\comparator/n2032 ) );
  inv \comparator/U2031  ( .a(\comparator/N14 ), .out(\comparator/n2031 ) );
  inv \comparator/U2030  ( .a(\comparator/N17 ), .out(\comparator/n2030 ) );
  inv \comparator/U2029  ( .a(\comparator/N16 ), .out(\comparator/n2029 ) );
  inv \comparator/U2028  ( .a(\comparator/N19 ), .out(\comparator/n2028 ) );
  inv \comparator/U2027  ( .a(\comparator/N18 ), .out(\comparator/n2027 ) );
  inv \comparator/U2026  ( .a(\comparator/N21 ), .out(\comparator/n2026 ) );
  inv \comparator/U2025  ( .a(\comparator/N20 ), .out(\comparator/n2025 ) );
  inv \comparator/U2024  ( .a(\comparator/N23 ), .out(\comparator/n2024 ) );
  inv \comparator/U2023  ( .a(\comparator/N22 ), .out(\comparator/n2023 ) );
  inv \comparator/U2022  ( .a(\comparator/N25 ), .out(\comparator/n2022 ) );
  inv \comparator/U2021  ( .a(\comparator/N24 ), .out(\comparator/n2021 ) );
  inv \comparator/U2020  ( .a(\comparator/N27 ), .out(\comparator/n2020 ) );
  inv \comparator/U2019  ( .a(\comparator/N26 ), .out(\comparator/n2019 ) );
  inv \comparator/U2018  ( .a(\comparator/N29 ), .out(\comparator/n2018 ) );
  inv \comparator/U2017  ( .a(\comparator/N28 ), .out(\comparator/n2017 ) );
  inv \comparator/U2016  ( .a(\comparator/N31 ), .out(\comparator/n2016 ) );
  inv \comparator/U2015  ( .a(\comparator/N30 ), .out(\comparator/n2015 ) );
  inv \comparator/U2014  ( .a(\comparator/N33 ), .out(\comparator/n2014 ) );
  inv \comparator/U2013  ( .a(\comparator/N32 ), .out(\comparator/n2013 ) );
  inv \comparator/U2012  ( .a(\comparator/N35 ), .out(\comparator/n2012 ) );
  inv \comparator/U2011  ( .a(\comparator/N34 ), .out(\comparator/n2011 ) );
  inv \comparator/U2010  ( .a(\comparator/N37 ), .out(\comparator/n2010 ) );
  inv \comparator/U2009  ( .a(\comparator/N36 ), .out(\comparator/n2009 ) );
  inv \comparator/U2008  ( .a(\comparator/N39 ), .out(\comparator/n2008 ) );
  inv \comparator/U2007  ( .a(\comparator/N38 ), .out(\comparator/n2007 ) );
  inv \comparator/U2006  ( .a(\comparator/N41 ), .out(\comparator/n2006 ) );
  inv \comparator/U2005  ( .a(\comparator/N40 ), .out(\comparator/n2005 ) );
  inv \comparator/U2004  ( .a(\comparator/N43 ), .out(\comparator/n2004 ) );
  inv \comparator/U2003  ( .a(\comparator/N42 ), .out(\comparator/n2003 ) );
  inv \comparator/U2002  ( .a(\comparator/N45 ), .out(\comparator/n2002 ) );
  inv \comparator/U2001  ( .a(\comparator/N44 ), .out(\comparator/n2001 ) );
  inv \comparator/U2000  ( .a(\comparator/N47 ), .out(\comparator/n2000 ) );
  inv \comparator/U1999  ( .a(\comparator/N46 ), .out(\comparator/n1999 ) );
  inv \comparator/U1998  ( .a(\comparator/N49 ), .out(\comparator/n1998 ) );
  inv \comparator/U1997  ( .a(\comparator/N48 ), .out(\comparator/n1997 ) );
  inv \comparator/U1996  ( .a(\comparator/N51 ), .out(\comparator/n1996 ) );
  inv \comparator/U1995  ( .a(\comparator/N50 ), .out(\comparator/n1995 ) );
  inv \comparator/U1994  ( .a(\comparator/N53 ), .out(\comparator/n1994 ) );
  inv \comparator/U1993  ( .a(\comparator/N52 ), .out(\comparator/n1993 ) );
  inv \comparator/U1992  ( .a(\comparator/N55 ), .out(\comparator/n1992 ) );
  inv \comparator/U1991  ( .a(\comparator/N54 ), .out(\comparator/n1991 ) );
  inv \comparator/U1990  ( .a(\comparator/N57 ), .out(\comparator/n1990 ) );
  inv \comparator/U1989  ( .a(\comparator/N56 ), .out(\comparator/n1989 ) );
  inv \comparator/U1988  ( .a(\comparator/N59 ), .out(\comparator/n1988 ) );
  inv \comparator/U1987  ( .a(\comparator/N58 ), .out(\comparator/n1987 ) );
  inv \comparator/U1986  ( .a(\comparator/N61 ), .out(\comparator/n1986 ) );
  inv \comparator/U1985  ( .a(\comparator/N60 ), .out(\comparator/n1985 ) );
  inv \comparator/U1984  ( .a(\comparator/N63 ), .out(\comparator/n1984 ) );
  inv \comparator/U1983  ( .a(\comparator/N62 ), .out(\comparator/n1983 ) );
  inv \comparator/U1982  ( .a(\comparator/N65 ), .out(\comparator/n1982 ) );
  inv \comparator/U1981  ( .a(\comparator/N64 ), .out(\comparator/n1981 ) );
  inv \comparator/U1980  ( .a(\comparator/N67 ), .out(\comparator/n1980 ) );
  inv \comparator/U1979  ( .a(\comparator/N66 ), .out(\comparator/n1979 ) );
  inv \comparator/U1978  ( .a(\comparator/N69 ), .out(\comparator/n1978 ) );
  inv \comparator/U1977  ( .a(\comparator/N68 ), .out(\comparator/n1977 ) );
  inv \comparator/U1976  ( .a(\comparator/N71 ), .out(\comparator/n1976 ) );
  inv \comparator/U1975  ( .a(\comparator/N70 ), .out(\comparator/n1975 ) );
  inv \comparator/U1974  ( .a(\comparator/N73 ), .out(\comparator/n1974 ) );
  inv \comparator/U1973  ( .a(\comparator/N72 ), .out(\comparator/n1973 ) );
  inv \comparator/U1972  ( .a(\comparator/N75 ), .out(\comparator/n1972 ) );
  inv \comparator/U1971  ( .a(\comparator/N74 ), .out(\comparator/n1971 ) );
  inv \comparator/U1970  ( .a(\comparator/N77 ), .out(\comparator/n1970 ) );
  inv \comparator/U1969  ( .a(\comparator/N76 ), .out(\comparator/n1969 ) );
  inv \comparator/U1968  ( .a(\comparator/N79 ), .out(\comparator/n1968 ) );
  inv \comparator/U1967  ( .a(\comparator/N78 ), .out(\comparator/n1967 ) );
  inv \comparator/U1966  ( .a(\comparator/N81 ), .out(\comparator/n1966 ) );
  inv \comparator/U1965  ( .a(\comparator/N80 ), .out(\comparator/n1965 ) );
  inv \comparator/U1964  ( .a(\comparator/N83 ), .out(\comparator/n1964 ) );
  inv \comparator/U1963  ( .a(\comparator/N82 ), .out(\comparator/n1963 ) );
  inv \comparator/U1962  ( .a(\comparator/N85 ), .out(\comparator/n1962 ) );
  inv \comparator/U1961  ( .a(\comparator/N84 ), .out(\comparator/n1961 ) );
  inv \comparator/U1960  ( .a(\comparator/N87 ), .out(\comparator/n1960 ) );
  inv \comparator/U1959  ( .a(\comparator/N86 ), .out(\comparator/n1959 ) );
  inv \comparator/U1958  ( .a(\comparator/N89 ), .out(\comparator/n1958 ) );
  inv \comparator/U1957  ( .a(\comparator/N88 ), .out(\comparator/n1957 ) );
  inv \comparator/U1956  ( .a(\comparator/N91 ), .out(\comparator/n1956 ) );
  inv \comparator/U1955  ( .a(\comparator/N90 ), .out(\comparator/n1955 ) );
  inv \comparator/U1954  ( .a(\comparator/N93 ), .out(\comparator/n1954 ) );
  inv \comparator/U1953  ( .a(\comparator/N92 ), .out(\comparator/n1953 ) );
  inv \comparator/U1952  ( .a(\comparator/N95 ), .out(\comparator/n1952 ) );
  inv \comparator/U1951  ( .a(\comparator/N94 ), .out(\comparator/n1951 ) );
  inv \comparator/U1950  ( .a(\comparator/N97 ), .out(\comparator/n1950 ) );
  inv \comparator/U1949  ( .a(\comparator/N96 ), .out(\comparator/n1949 ) );
  inv \comparator/U1948  ( .a(\comparator/N99 ), .out(\comparator/n1948 ) );
  inv \comparator/U1947  ( .a(\comparator/N98 ), .out(\comparator/n1947 ) );
  inv \comparator/U1946  ( .a(\comparator/N101 ), .out(\comparator/n1946 ) );
  inv \comparator/U1945  ( .a(\comparator/N100 ), .out(\comparator/n1945 ) );
  inv \comparator/U1944  ( .a(\comparator/N103 ), .out(\comparator/n1944 ) );
  inv \comparator/U1943  ( .a(\comparator/N102 ), .out(\comparator/n1943 ) );
  inv \comparator/U1942  ( .a(\comparator/N105 ), .out(\comparator/n1942 ) );
  inv \comparator/U1941  ( .a(\comparator/N104 ), .out(\comparator/n1941 ) );
  inv \comparator/U1940  ( .a(\comparator/N107 ), .out(\comparator/n1940 ) );
  inv \comparator/U1939  ( .a(\comparator/N106 ), .out(\comparator/n1939 ) );
  inv \comparator/U1938  ( .a(\comparator/N109 ), .out(\comparator/n1938 ) );
  inv \comparator/U1937  ( .a(\comparator/N108 ), .out(\comparator/n1937 ) );
  inv \comparator/U1936  ( .a(\comparator/N111 ), .out(\comparator/n1936 ) );
  inv \comparator/U1935  ( .a(\comparator/N110 ), .out(\comparator/n1935 ) );
  inv \comparator/U1934  ( .a(\comparator/N113 ), .out(\comparator/n1934 ) );
  inv \comparator/U1933  ( .a(\comparator/N112 ), .out(\comparator/n1933 ) );
  inv \comparator/U1932  ( .a(\comparator/N115 ), .out(\comparator/n1932 ) );
  inv \comparator/U1931  ( .a(\comparator/N114 ), .out(\comparator/n1931 ) );
  inv \comparator/U1930  ( .a(\comparator/N117 ), .out(\comparator/n1930 ) );
  inv \comparator/U1929  ( .a(\comparator/N116 ), .out(\comparator/n1929 ) );
  inv \comparator/U1928  ( .a(\comparator/N119 ), .out(\comparator/n1928 ) );
  inv \comparator/U1927  ( .a(\comparator/N118 ), .out(\comparator/n1927 ) );
  inv \comparator/U1926  ( .a(\comparator/N121 ), .out(\comparator/n1926 ) );
  inv \comparator/U1925  ( .a(\comparator/N120 ), .out(\comparator/n1925 ) );
  inv \comparator/U1924  ( .a(\comparator/N123 ), .out(\comparator/n1924 ) );
  inv \comparator/U1923  ( .a(\comparator/N122 ), .out(\comparator/n1923 ) );
  inv \comparator/U1922  ( .a(\comparator/N125 ), .out(\comparator/n1922 ) );
  inv \comparator/U1921  ( .a(\comparator/N124 ), .out(\comparator/n1921 ) );
  inv \comparator/U1920  ( .a(\comparator/N127 ), .out(\comparator/n1920 ) );
  inv \comparator/U1919  ( .a(\comparator/N126 ), .out(\comparator/n1919 ) );
  inv \comparator/U1918  ( .a(\comparator/N129 ), .out(\comparator/n1918 ) );
  inv \comparator/U1917  ( .a(\comparator/N128 ), .out(\comparator/n1917 ) );
  inv \comparator/U1916  ( .a(\comparator/N131 ), .out(\comparator/n1916 ) );
  inv \comparator/U1915  ( .a(\comparator/N130 ), .out(\comparator/n1915 ) );
  inv \comparator/U1914  ( .a(\comparator/N133 ), .out(\comparator/n1914 ) );
  inv \comparator/U1913  ( .a(\comparator/N132 ), .out(\comparator/n1913 ) );
  inv \comparator/U1912  ( .a(\comparator/N135 ), .out(\comparator/n1912 ) );
  inv \comparator/U1911  ( .a(\comparator/N134 ), .out(\comparator/n1911 ) );
  inv \comparator/U1910  ( .a(\comparator/N137 ), .out(\comparator/n1910 ) );
  inv \comparator/U1909  ( .a(\comparator/N136 ), .out(\comparator/n1909 ) );
  inv \comparator/U1908  ( .a(\comparator/N139 ), .out(\comparator/n1908 ) );
  inv \comparator/U1907  ( .a(\comparator/N138 ), .out(\comparator/n1907 ) );
  inv \comparator/U1906  ( .a(\comparator/N141 ), .out(\comparator/n1906 ) );
  inv \comparator/U1905  ( .a(\comparator/N140 ), .out(\comparator/n1905 ) );
  inv \comparator/U1904  ( .a(\comparator/N143 ), .out(\comparator/n1904 ) );
  inv \comparator/U1903  ( .a(\comparator/N142 ), .out(\comparator/n1903 ) );
  inv \comparator/U1902  ( .a(\comparator/N145 ), .out(\comparator/n1902 ) );
  inv \comparator/U1901  ( .a(\comparator/N144 ), .out(\comparator/n1901 ) );
  inv \comparator/U1900  ( .a(\comparator/N147 ), .out(\comparator/n1900 ) );
  inv \comparator/U1899  ( .a(\comparator/N146 ), .out(\comparator/n1899 ) );
  inv \comparator/U1898  ( .a(\comparator/N149 ), .out(\comparator/n1898 ) );
  inv \comparator/U1897  ( .a(\comparator/N148 ), .out(\comparator/n1897 ) );
  inv \comparator/U1896  ( .a(\comparator/N151 ), .out(\comparator/n1896 ) );
  inv \comparator/U1895  ( .a(\comparator/N150 ), .out(\comparator/n1895 ) );
  inv \comparator/U1894  ( .a(\comparator/N153 ), .out(\comparator/n1894 ) );
  inv \comparator/U1893  ( .a(\comparator/N152 ), .out(\comparator/n1893 ) );
  inv \comparator/U1892  ( .a(\comparator/N155 ), .out(\comparator/n1892 ) );
  inv \comparator/U1891  ( .a(\comparator/N154 ), .out(\comparator/n1891 ) );
  inv \comparator/U1890  ( .a(\comparator/N157 ), .out(\comparator/n1890 ) );
  inv \comparator/U1889  ( .a(\comparator/N156 ), .out(\comparator/n1889 ) );
  inv \comparator/U1888  ( .a(\comparator/N159 ), .out(\comparator/n1888 ) );
  inv \comparator/U1887  ( .a(\comparator/N158 ), .out(\comparator/n1887 ) );
  inv \comparator/U1886  ( .a(\comparator/N161 ), .out(\comparator/n1886 ) );
  inv \comparator/U1885  ( .a(\comparator/N160 ), .out(\comparator/n1885 ) );
  inv \comparator/U1884  ( .a(\comparator/N163 ), .out(\comparator/n1884 ) );
  inv \comparator/U1883  ( .a(\comparator/N162 ), .out(\comparator/n1883 ) );
  inv \comparator/U1882  ( .a(\comparator/N165 ), .out(\comparator/n1882 ) );
  inv \comparator/U1881  ( .a(\comparator/N164 ), .out(\comparator/n1881 ) );
  inv \comparator/U1880  ( .a(\comparator/N167 ), .out(\comparator/n1880 ) );
  inv \comparator/U1879  ( .a(\comparator/N166 ), .out(\comparator/n1879 ) );
  inv \comparator/U1878  ( .a(\comparator/N169 ), .out(\comparator/n1878 ) );
  inv \comparator/U1877  ( .a(\comparator/N168 ), .out(\comparator/n1877 ) );
  inv \comparator/U1876  ( .a(\comparator/N171 ), .out(\comparator/n1876 ) );
  inv \comparator/U1875  ( .a(\comparator/N170 ), .out(\comparator/n1875 ) );
  inv \comparator/U1874  ( .a(\comparator/N173 ), .out(\comparator/n1874 ) );
  inv \comparator/U1873  ( .a(\comparator/N172 ), .out(\comparator/n1873 ) );
  inv \comparator/U1872  ( .a(\comparator/N175 ), .out(\comparator/n1872 ) );
  inv \comparator/U1871  ( .a(\comparator/N174 ), .out(\comparator/n1871 ) );
  inv \comparator/U1870  ( .a(\comparator/N177 ), .out(\comparator/n1870 ) );
  inv \comparator/U1869  ( .a(\comparator/N176 ), .out(\comparator/n1869 ) );
  inv \comparator/U1868  ( .a(\comparator/N179 ), .out(\comparator/n1868 ) );
  inv \comparator/U1867  ( .a(\comparator/N178 ), .out(\comparator/n1867 ) );
  inv \comparator/U1866  ( .a(\comparator/N181 ), .out(\comparator/n1866 ) );
  inv \comparator/U1865  ( .a(\comparator/N180 ), .out(\comparator/n1865 ) );
  inv \comparator/U1864  ( .a(\comparator/N183 ), .out(\comparator/n1864 ) );
  inv \comparator/U1863  ( .a(\comparator/N182 ), .out(\comparator/n1863 ) );
  inv \comparator/U1862  ( .a(\comparator/N185 ), .out(\comparator/n1862 ) );
  inv \comparator/U1861  ( .a(\comparator/N184 ), .out(\comparator/n1861 ) );
  inv \comparator/U1860  ( .a(\comparator/N187 ), .out(\comparator/n1860 ) );
  inv \comparator/U1859  ( .a(\comparator/N186 ), .out(\comparator/n1859 ) );
  inv \comparator/U1858  ( .a(\comparator/N189 ), .out(\comparator/n1858 ) );
  inv \comparator/U1857  ( .a(\comparator/N188 ), .out(\comparator/n1857 ) );
  inv \comparator/U1856  ( .a(\comparator/N191 ), .out(\comparator/n1856 ) );
  inv \comparator/U1855  ( .a(\comparator/N190 ), .out(\comparator/n1855 ) );
  inv \comparator/U1854  ( .a(\comparator/N193 ), .out(\comparator/n1854 ) );
  inv \comparator/U1853  ( .a(\comparator/N192 ), .out(\comparator/n1853 ) );
  inv \comparator/U1852  ( .a(\comparator/N195 ), .out(\comparator/n1852 ) );
  inv \comparator/U1851  ( .a(\comparator/N194 ), .out(\comparator/n1851 ) );
  inv \comparator/U1850  ( .a(\comparator/N197 ), .out(\comparator/n1850 ) );
  inv \comparator/U1849  ( .a(\comparator/N196 ), .out(\comparator/n1849 ) );
  inv \comparator/U1848  ( .a(\comparator/N199 ), .out(\comparator/n1848 ) );
  inv \comparator/U1847  ( .a(\comparator/N198 ), .out(\comparator/n1847 ) );
  inv \comparator/U1846  ( .a(\comparator/N201 ), .out(\comparator/n1846 ) );
  inv \comparator/U1845  ( .a(\comparator/N200 ), .out(\comparator/n1845 ) );
  inv \comparator/U1844  ( .a(\comparator/N203 ), .out(\comparator/n1844 ) );
  inv \comparator/U1843  ( .a(\comparator/N202 ), .out(\comparator/n1843 ) );
  inv \comparator/U1842  ( .a(\comparator/N205 ), .out(\comparator/n1842 ) );
  inv \comparator/U1841  ( .a(\comparator/N204 ), .out(\comparator/n1841 ) );
  inv \comparator/U1840  ( .a(\comparator/N207 ), .out(\comparator/n1840 ) );
  inv \comparator/U1839  ( .a(\comparator/N206 ), .out(\comparator/n1839 ) );
  inv \comparator/U1838  ( .a(\comparator/N209 ), .out(\comparator/n1838 ) );
  inv \comparator/U1837  ( .a(\comparator/N208 ), .out(\comparator/n1837 ) );
  inv \comparator/U1836  ( .a(\comparator/N211 ), .out(\comparator/n1836 ) );
  inv \comparator/U1835  ( .a(\comparator/N210 ), .out(\comparator/n1835 ) );
  inv \comparator/U1834  ( .a(\comparator/N213 ), .out(\comparator/n1834 ) );
  inv \comparator/U1833  ( .a(\comparator/N212 ), .out(\comparator/n1833 ) );
  inv \comparator/U1832  ( .a(\comparator/N215 ), .out(\comparator/n1832 ) );
  inv \comparator/U1831  ( .a(\comparator/N214 ), .out(\comparator/n1831 ) );
  inv \comparator/U1830  ( .a(\comparator/N217 ), .out(\comparator/n1830 ) );
  inv \comparator/U1829  ( .a(\comparator/N216 ), .out(\comparator/n1829 ) );
  inv \comparator/U1828  ( .a(\comparator/N219 ), .out(\comparator/n1828 ) );
  inv \comparator/U1827  ( .a(\comparator/N218 ), .out(\comparator/n1827 ) );
  inv \comparator/U1826  ( .a(\comparator/N221 ), .out(\comparator/n1826 ) );
  inv \comparator/U1825  ( .a(\comparator/N220 ), .out(\comparator/n1825 ) );
  inv \comparator/U1824  ( .a(\comparator/N223 ), .out(\comparator/n1824 ) );
  inv \comparator/U1823  ( .a(\comparator/N222 ), .out(\comparator/n1823 ) );
  inv \comparator/U1822  ( .a(\comparator/N225 ), .out(\comparator/n1822 ) );
  inv \comparator/U1821  ( .a(\comparator/N224 ), .out(\comparator/n1821 ) );
  inv \comparator/U1820  ( .a(\comparator/N227 ), .out(\comparator/n1820 ) );
  inv \comparator/U1819  ( .a(\comparator/N226 ), .out(\comparator/n1819 ) );
  inv \comparator/U1818  ( .a(\comparator/N229 ), .out(\comparator/n1818 ) );
  inv \comparator/U1817  ( .a(\comparator/N228 ), .out(\comparator/n1817 ) );
  inv \comparator/U1816  ( .a(\comparator/N231 ), .out(\comparator/n1816 ) );
  inv \comparator/U1815  ( .a(\comparator/N230 ), .out(\comparator/n1815 ) );
  inv \comparator/U1814  ( .a(\comparator/N233 ), .out(\comparator/n1814 ) );
  inv \comparator/U1813  ( .a(\comparator/N232 ), .out(\comparator/n1813 ) );
  inv \comparator/U1812  ( .a(\comparator/N235 ), .out(\comparator/n1812 ) );
  inv \comparator/U1811  ( .a(\comparator/N234 ), .out(\comparator/n1811 ) );
  inv \comparator/U1810  ( .a(\comparator/N237 ), .out(\comparator/n1810 ) );
  inv \comparator/U1809  ( .a(\comparator/N236 ), .out(\comparator/n1809 ) );
  inv \comparator/U1808  ( .a(\comparator/N239 ), .out(\comparator/n1808 ) );
  inv \comparator/U1807  ( .a(\comparator/N238 ), .out(\comparator/n1807 ) );
  inv \comparator/U1806  ( .a(\comparator/N241 ), .out(\comparator/n1806 ) );
  inv \comparator/U1805  ( .a(\comparator/N240 ), .out(\comparator/n1805 ) );
  inv \comparator/U1804  ( .a(\comparator/N243 ), .out(\comparator/n1804 ) );
  inv \comparator/U1803  ( .a(\comparator/N242 ), .out(\comparator/n1803 ) );
  inv \comparator/U1802  ( .a(\comparator/N245 ), .out(\comparator/n1802 ) );
  inv \comparator/U1801  ( .a(\comparator/N244 ), .out(\comparator/n1801 ) );
  inv \comparator/U1800  ( .a(\comparator/N247 ), .out(\comparator/n1800 ) );
  inv \comparator/U1799  ( .a(\comparator/N246 ), .out(\comparator/n1799 ) );
  inv \comparator/U1798  ( .a(\comparator/N249 ), .out(\comparator/n1798 ) );
  inv \comparator/U1797  ( .a(\comparator/N248 ), .out(\comparator/n1797 ) );
  inv \comparator/U1796  ( .a(\comparator/N251 ), .out(\comparator/n1796 ) );
  inv \comparator/U1795  ( .a(\comparator/N250 ), .out(\comparator/n1795 ) );
  inv \comparator/U1794  ( .a(\comparator/N253 ), .out(\comparator/n1794 ) );
  inv \comparator/U1793  ( .a(\comparator/N252 ), .out(\comparator/n1793 ) );
  inv \comparator/U1792  ( .a(\comparator/N255 ), .out(\comparator/n1792 ) );
  inv \comparator/U1791  ( .a(\comparator/N254 ), .out(\comparator/n1791 ) );
  inv \comparator/U1790  ( .a(\comparator/N257 ), .out(\comparator/n1790 ) );
  inv \comparator/U1789  ( .a(\comparator/N256 ), .out(\comparator/n1789 ) );
  inv \comparator/U1788  ( .a(\comparator/N259 ), .out(\comparator/n1788 ) );
  inv \comparator/U1787  ( .a(\comparator/N258 ), .out(\comparator/n1787 ) );
  inv \comparator/U1786  ( .a(\comparator/N261 ), .out(\comparator/n1786 ) );
  inv \comparator/U1785  ( .a(\comparator/N260 ), .out(\comparator/n1785 ) );
  inv \comparator/U1784  ( .a(\comparator/N263 ), .out(\comparator/n1784 ) );
  inv \comparator/U1783  ( .a(\comparator/N262 ), .out(\comparator/n1783 ) );
  inv \comparator/U1782  ( .a(\comparator/N265 ), .out(\comparator/n1782 ) );
  inv \comparator/U1781  ( .a(\comparator/N264 ), .out(\comparator/n1781 ) );
  inv \comparator/U1780  ( .a(\comparator/N267 ), .out(\comparator/n1780 ) );
  inv \comparator/U1779  ( .a(\comparator/N266 ), .out(\comparator/n1779 ) );
  inv \comparator/U1778  ( .a(\comparator/N269 ), .out(\comparator/n1778 ) );
  inv \comparator/U1777  ( .a(\comparator/N268 ), .out(\comparator/n1777 ) );
  inv \comparator/U1776  ( .a(\comparator/N271 ), .out(\comparator/n1776 ) );
  inv \comparator/U1775  ( .a(\comparator/N270 ), .out(\comparator/n1775 ) );
  inv \comparator/U1774  ( .a(\comparator/N273 ), .out(\comparator/n1774 ) );
  inv \comparator/U1773  ( .a(\comparator/N272 ), .out(\comparator/n1773 ) );
  inv \comparator/U1772  ( .a(\comparator/N275 ), .out(\comparator/n1772 ) );
  inv \comparator/U1771  ( .a(\comparator/N274 ), .out(\comparator/n1771 ) );
  inv \comparator/U1770  ( .a(\comparator/N277 ), .out(\comparator/n1770 ) );
  inv \comparator/U1769  ( .a(\comparator/N276 ), .out(\comparator/n1769 ) );
  inv \comparator/U1768  ( .a(\comparator/N279 ), .out(\comparator/n1768 ) );
  inv \comparator/U1767  ( .a(\comparator/N278 ), .out(\comparator/n1767 ) );
  inv \comparator/U1766  ( .a(\comparator/N281 ), .out(\comparator/n1766 ) );
  inv \comparator/U1765  ( .a(\comparator/N280 ), .out(\comparator/n1765 ) );
  inv \comparator/U1764  ( .a(\comparator/N283 ), .out(\comparator/n1764 ) );
  inv \comparator/U1763  ( .a(\comparator/N282 ), .out(\comparator/n1763 ) );
  inv \comparator/U1762  ( .a(\comparator/N285 ), .out(\comparator/n1762 ) );
  inv \comparator/U1761  ( .a(\comparator/N284 ), .out(\comparator/n1761 ) );
  inv \comparator/U1760  ( .a(\comparator/N287 ), .out(\comparator/n1760 ) );
  inv \comparator/U1759  ( .a(\comparator/N286 ), .out(\comparator/n1759 ) );
  inv \comparator/U1758  ( .a(\comparator/N289 ), .out(\comparator/n1758 ) );
  inv \comparator/U1757  ( .a(\comparator/N288 ), .out(\comparator/n1757 ) );
  inv \comparator/U1756  ( .a(\comparator/N291 ), .out(\comparator/n1756 ) );
  inv \comparator/U1755  ( .a(\comparator/N290 ), .out(\comparator/n1755 ) );
  inv \comparator/U1754  ( .a(\comparator/N293 ), .out(\comparator/n1754 ) );
  inv \comparator/U1753  ( .a(\comparator/N292 ), .out(\comparator/n1753 ) );
  inv \comparator/U1752  ( .a(\comparator/N295 ), .out(\comparator/n1752 ) );
  inv \comparator/U1751  ( .a(\comparator/N294 ), .out(\comparator/n1751 ) );
  inv \comparator/U1750  ( .a(\comparator/N297 ), .out(\comparator/n1750 ) );
  inv \comparator/U1749  ( .a(\comparator/N296 ), .out(\comparator/n1749 ) );
  inv \comparator/U1748  ( .a(\comparator/N299 ), .out(\comparator/n1748 ) );
  inv \comparator/U1747  ( .a(\comparator/N298 ), .out(\comparator/n1747 ) );
  inv \comparator/U1746  ( .a(\comparator/N301 ), .out(\comparator/n1746 ) );
  inv \comparator/U1745  ( .a(\comparator/N300 ), .out(\comparator/n1745 ) );
  inv \comparator/U1744  ( .a(\comparator/N303 ), .out(\comparator/n1744 ) );
  inv \comparator/U1743  ( .a(\comparator/N302 ), .out(\comparator/n1743 ) );
  inv \comparator/U1742  ( .a(\comparator/N305 ), .out(\comparator/n1742 ) );
  inv \comparator/U1741  ( .a(\comparator/N304 ), .out(\comparator/n1741 ) );
  inv \comparator/U1740  ( .a(\comparator/N307 ), .out(\comparator/n1740 ) );
  inv \comparator/U1739  ( .a(\comparator/N306 ), .out(\comparator/n1739 ) );
  inv \comparator/U1738  ( .a(\comparator/N309 ), .out(\comparator/n1738 ) );
  inv \comparator/U1737  ( .a(\comparator/N308 ), .out(\comparator/n1737 ) );
  inv \comparator/U1736  ( .a(\comparator/N311 ), .out(\comparator/n1736 ) );
  inv \comparator/U1735  ( .a(\comparator/N310 ), .out(\comparator/n1735 ) );
  inv \comparator/U1734  ( .a(\comparator/N313 ), .out(\comparator/n1734 ) );
  inv \comparator/U1733  ( .a(\comparator/N312 ), .out(\comparator/n1733 ) );
  inv \comparator/U1732  ( .a(\comparator/N315 ), .out(\comparator/n1732 ) );
  inv \comparator/U1731  ( .a(\comparator/N314 ), .out(\comparator/n1731 ) );
  inv \comparator/U1730  ( .a(\comparator/N317 ), .out(\comparator/n1730 ) );
  inv \comparator/U1729  ( .a(\comparator/N316 ), .out(\comparator/n1729 ) );
  inv \comparator/U1728  ( .a(\comparator/N319 ), .out(\comparator/n1728 ) );
  inv \comparator/U1727  ( .a(\comparator/N318 ), .out(\comparator/n1727 ) );
  inv \comparator/U1726  ( .a(\comparator/N321 ), .out(\comparator/n1726 ) );
  inv \comparator/U1725  ( .a(\comparator/N320 ), .out(\comparator/n1725 ) );
  inv \comparator/U1724  ( .a(\comparator/N323 ), .out(\comparator/n1724 ) );
  inv \comparator/U1723  ( .a(\comparator/N322 ), .out(\comparator/n1723 ) );
  inv \comparator/U1722  ( .a(\comparator/N325 ), .out(\comparator/n1722 ) );
  inv \comparator/U1721  ( .a(\comparator/N324 ), .out(\comparator/n1721 ) );
  inv \comparator/U1720  ( .a(\comparator/N327 ), .out(\comparator/n1720 ) );
  inv \comparator/U1719  ( .a(\comparator/N326 ), .out(\comparator/n1719 ) );
  inv \comparator/U1718  ( .a(\comparator/N329 ), .out(\comparator/n1718 ) );
  inv \comparator/U1717  ( .a(\comparator/N328 ), .out(\comparator/n1717 ) );
  inv \comparator/U1716  ( .a(\comparator/N331 ), .out(\comparator/n1716 ) );
  inv \comparator/U1715  ( .a(\comparator/N330 ), .out(\comparator/n1715 ) );
  inv \comparator/U1714  ( .a(\comparator/N333 ), .out(\comparator/n1714 ) );
  inv \comparator/U1713  ( .a(\comparator/N332 ), .out(\comparator/n1713 ) );
  inv \comparator/U1712  ( .a(\comparator/N335 ), .out(\comparator/n1712 ) );
  inv \comparator/U1711  ( .a(\comparator/N334 ), .out(\comparator/n1711 ) );
  inv \comparator/U1710  ( .a(\comparator/N337 ), .out(\comparator/n1710 ) );
  inv \comparator/U1709  ( .a(\comparator/N336 ), .out(\comparator/n1709 ) );
  inv \comparator/U1708  ( .a(\comparator/N339 ), .out(\comparator/n1708 ) );
  inv \comparator/U1707  ( .a(\comparator/N338 ), .out(\comparator/n1707 ) );
  inv \comparator/U1706  ( .a(\comparator/N341 ), .out(\comparator/n1706 ) );
  inv \comparator/U1705  ( .a(\comparator/N340 ), .out(\comparator/n1705 ) );
  inv \comparator/U1704  ( .a(\comparator/N343 ), .out(\comparator/n1704 ) );
  inv \comparator/U1703  ( .a(\comparator/N342 ), .out(\comparator/n1703 ) );
  inv \comparator/U1702  ( .a(\comparator/N345 ), .out(\comparator/n1702 ) );
  inv \comparator/U1701  ( .a(\comparator/N344 ), .out(\comparator/n1701 ) );
  inv \comparator/U1700  ( .a(\comparator/N347 ), .out(\comparator/n1700 ) );
  inv \comparator/U1699  ( .a(\comparator/N346 ), .out(\comparator/n1699 ) );
  inv \comparator/U1698  ( .a(\comparator/N349 ), .out(\comparator/n1698 ) );
  inv \comparator/U1697  ( .a(\comparator/N348 ), .out(\comparator/n1697 ) );
  inv \comparator/U1696  ( .a(\comparator/N351 ), .out(\comparator/n1696 ) );
  inv \comparator/U1695  ( .a(\comparator/N350 ), .out(\comparator/n1695 ) );
  inv \comparator/U1694  ( .a(\comparator/N353 ), .out(\comparator/n1694 ) );
  inv \comparator/U1693  ( .a(\comparator/N352 ), .out(\comparator/n1693 ) );
  inv \comparator/U1692  ( .a(\comparator/N355 ), .out(\comparator/n1692 ) );
  inv \comparator/U1691  ( .a(\comparator/N354 ), .out(\comparator/n1691 ) );
  inv \comparator/U1690  ( .a(\comparator/N357 ), .out(\comparator/n1690 ) );
  inv \comparator/U1689  ( .a(\comparator/N356 ), .out(\comparator/n1689 ) );
  inv \comparator/U1688  ( .a(\comparator/N359 ), .out(\comparator/n1688 ) );
  inv \comparator/U1687  ( .a(\comparator/N358 ), .out(\comparator/n1687 ) );
  inv \comparator/U1686  ( .a(\comparator/N361 ), .out(\comparator/n1686 ) );
  inv \comparator/U1685  ( .a(\comparator/N360 ), .out(\comparator/n1685 ) );
  inv \comparator/U1684  ( .a(\comparator/N363 ), .out(\comparator/n1684 ) );
  inv \comparator/U1683  ( .a(\comparator/N362 ), .out(\comparator/n1683 ) );
  inv \comparator/U1682  ( .a(\comparator/N365 ), .out(\comparator/n1682 ) );
  inv \comparator/U1681  ( .a(\comparator/N364 ), .out(\comparator/n1681 ) );
  inv \comparator/U1680  ( .a(\comparator/N367 ), .out(\comparator/n1680 ) );
  inv \comparator/U1679  ( .a(\comparator/N366 ), .out(\comparator/n1679 ) );
  inv \comparator/U1678  ( .a(\comparator/N369 ), .out(\comparator/n1678 ) );
  inv \comparator/U1677  ( .a(\comparator/N368 ), .out(\comparator/n1677 ) );
  inv \comparator/U1676  ( .a(\comparator/N371 ), .out(\comparator/n1676 ) );
  inv \comparator/U1675  ( .a(\comparator/N370 ), .out(\comparator/n1675 ) );
  inv \comparator/U1674  ( .a(\comparator/N373 ), .out(\comparator/n1674 ) );
  inv \comparator/U1673  ( .a(\comparator/N372 ), .out(\comparator/n1673 ) );
  inv \comparator/U1672  ( .a(\comparator/N375 ), .out(\comparator/n1672 ) );
  inv \comparator/U1671  ( .a(\comparator/N374 ), .out(\comparator/n1671 ) );
  inv \comparator/U1670  ( .a(\comparator/N377 ), .out(\comparator/n1670 ) );
  inv \comparator/U1669  ( .a(\comparator/N376 ), .out(\comparator/n1669 ) );
  inv \comparator/U1668  ( .a(\comparator/N379 ), .out(\comparator/n1668 ) );
  inv \comparator/U1667  ( .a(\comparator/N378 ), .out(\comparator/n1667 ) );
  inv \comparator/U1666  ( .a(\comparator/N381 ), .out(\comparator/n1666 ) );
  inv \comparator/U1665  ( .a(\comparator/N380 ), .out(\comparator/n1665 ) );
  inv \comparator/U1664  ( .a(\comparator/N383 ), .out(\comparator/n1664 ) );
  inv \comparator/U1663  ( .a(\comparator/N382 ), .out(\comparator/n1663 ) );
  inv \comparator/U1662  ( .a(\comparator/N385 ), .out(\comparator/n1662 ) );
  inv \comparator/U1661  ( .a(\comparator/N384 ), .out(\comparator/n1661 ) );
  inv \comparator/U1660  ( .a(\comparator/N387 ), .out(\comparator/n1660 ) );
  inv \comparator/U1659  ( .a(\comparator/N386 ), .out(\comparator/n1659 ) );
  inv \comparator/U1658  ( .a(\comparator/N389 ), .out(\comparator/n1658 ) );
  inv \comparator/U1657  ( .a(\comparator/N388 ), .out(\comparator/n1657 ) );
  inv \comparator/U1656  ( .a(\comparator/N391 ), .out(\comparator/n1656 ) );
  inv \comparator/U1655  ( .a(\comparator/N390 ), .out(\comparator/n1655 ) );
  inv \comparator/U1654  ( .a(\comparator/N393 ), .out(\comparator/n1654 ) );
  inv \comparator/U1653  ( .a(\comparator/N392 ), .out(\comparator/n1653 ) );
  inv \comparator/U1652  ( .a(\comparator/N395 ), .out(\comparator/n1652 ) );
  inv \comparator/U1651  ( .a(\comparator/N394 ), .out(\comparator/n1651 ) );
  inv \comparator/U1650  ( .a(\comparator/N397 ), .out(\comparator/n1650 ) );
  inv \comparator/U1649  ( .a(\comparator/N396 ), .out(\comparator/n1649 ) );
  inv \comparator/U1648  ( .a(\comparator/N399 ), .out(\comparator/n1648 ) );
  inv \comparator/U1647  ( .a(\comparator/N398 ), .out(\comparator/n1647 ) );
  inv \comparator/U1646  ( .a(\comparator/N401 ), .out(\comparator/n1646 ) );
  inv \comparator/U1645  ( .a(\comparator/N400 ), .out(\comparator/n1645 ) );
  inv \comparator/U1644  ( .a(\comparator/N403 ), .out(\comparator/n1644 ) );
  inv \comparator/U1643  ( .a(\comparator/N402 ), .out(\comparator/n1643 ) );
  inv \comparator/U1642  ( .a(\comparator/N405 ), .out(\comparator/n1642 ) );
  inv \comparator/U1641  ( .a(\comparator/N404 ), .out(\comparator/n1641 ) );
  inv \comparator/U1640  ( .a(\comparator/N407 ), .out(\comparator/n1640 ) );
  inv \comparator/U1639  ( .a(\comparator/N406 ), .out(\comparator/n1639 ) );
  inv \comparator/U1638  ( .a(\comparator/N409 ), .out(\comparator/n1638 ) );
  inv \comparator/U1637  ( .a(\comparator/N408 ), .out(\comparator/n1637 ) );
  inv \comparator/U1636  ( .a(\comparator/N411 ), .out(\comparator/n1636 ) );
  inv \comparator/U1635  ( .a(\comparator/N410 ), .out(\comparator/n1635 ) );
  inv \comparator/U1634  ( .a(\comparator/N413 ), .out(\comparator/n1634 ) );
  inv \comparator/U1633  ( .a(\comparator/N412 ), .out(\comparator/n1633 ) );
  inv \comparator/U1632  ( .a(\comparator/N415 ), .out(\comparator/n1632 ) );
  inv \comparator/U1631  ( .a(\comparator/N414 ), .out(\comparator/n1631 ) );
  inv \comparator/U1630  ( .a(\comparator/N417 ), .out(\comparator/n1630 ) );
  inv \comparator/U1629  ( .a(\comparator/N416 ), .out(\comparator/n1629 ) );
  inv \comparator/U1628  ( .a(\comparator/N419 ), .out(\comparator/n1628 ) );
  inv \comparator/U1627  ( .a(\comparator/N418 ), .out(\comparator/n1627 ) );
  inv \comparator/U1626  ( .a(\comparator/N421 ), .out(\comparator/n1626 ) );
  inv \comparator/U1625  ( .a(\comparator/N420 ), .out(\comparator/n1625 ) );
  inv \comparator/U1624  ( .a(\comparator/N423 ), .out(\comparator/n1624 ) );
  inv \comparator/U1623  ( .a(\comparator/N422 ), .out(\comparator/n1623 ) );
  inv \comparator/U1622  ( .a(\comparator/N425 ), .out(\comparator/n1622 ) );
  inv \comparator/U1621  ( .a(\comparator/N424 ), .out(\comparator/n1621 ) );
  inv \comparator/U1620  ( .a(\comparator/N427 ), .out(\comparator/n1620 ) );
  inv \comparator/U1619  ( .a(\comparator/N426 ), .out(\comparator/n1619 ) );
  inv \comparator/U1618  ( .a(\comparator/N429 ), .out(\comparator/n1618 ) );
  inv \comparator/U1617  ( .a(\comparator/N428 ), .out(\comparator/n1617 ) );
  inv \comparator/U1616  ( .a(\comparator/N431 ), .out(\comparator/n1616 ) );
  inv \comparator/U1615  ( .a(\comparator/N430 ), .out(\comparator/n1615 ) );
  inv \comparator/U1614  ( .a(\comparator/N433 ), .out(\comparator/n1614 ) );
  inv \comparator/U1613  ( .a(\comparator/N432 ), .out(\comparator/n1613 ) );
  inv \comparator/U1612  ( .a(\comparator/N435 ), .out(\comparator/n1612 ) );
  inv \comparator/U1611  ( .a(\comparator/N434 ), .out(\comparator/n1611 ) );
  inv \comparator/U1610  ( .a(\comparator/N437 ), .out(\comparator/n1610 ) );
  inv \comparator/U1609  ( .a(\comparator/N436 ), .out(\comparator/n1609 ) );
  inv \comparator/U1608  ( .a(\comparator/N439 ), .out(\comparator/n1608 ) );
  inv \comparator/U1607  ( .a(\comparator/N438 ), .out(\comparator/n1607 ) );
  inv \comparator/U1606  ( .a(\comparator/N441 ), .out(\comparator/n1606 ) );
  inv \comparator/U1605  ( .a(\comparator/N440 ), .out(\comparator/n1605 ) );
  inv \comparator/U1604  ( .a(\comparator/N443 ), .out(\comparator/n1604 ) );
  inv \comparator/U1603  ( .a(\comparator/N442 ), .out(\comparator/n1603 ) );
  inv \comparator/U1602  ( .a(\comparator/N445 ), .out(\comparator/n1602 ) );
  inv \comparator/U1601  ( .a(\comparator/N444 ), .out(\comparator/n1601 ) );
  inv \comparator/U1600  ( .a(\comparator/N447 ), .out(\comparator/n1600 ) );
  inv \comparator/U1599  ( .a(\comparator/N446 ), .out(\comparator/n1599 ) );
  inv \comparator/U1598  ( .a(\comparator/N449 ), .out(\comparator/n1598 ) );
  inv \comparator/U1597  ( .a(\comparator/N448 ), .out(\comparator/n1597 ) );
  inv \comparator/U1596  ( .a(\comparator/N451 ), .out(\comparator/n1596 ) );
  inv \comparator/U1595  ( .a(\comparator/N450 ), .out(\comparator/n1595 ) );
  inv \comparator/U1594  ( .a(\comparator/N453 ), .out(\comparator/n1594 ) );
  inv \comparator/U1593  ( .a(\comparator/N452 ), .out(\comparator/n1593 ) );
  inv \comparator/U1592  ( .a(\comparator/N455 ), .out(\comparator/n1592 ) );
  inv \comparator/U1591  ( .a(\comparator/N454 ), .out(\comparator/n1591 ) );
  inv \comparator/U1590  ( .a(\comparator/N457 ), .out(\comparator/n1590 ) );
  inv \comparator/U1589  ( .a(\comparator/N456 ), .out(\comparator/n1589 ) );
  inv \comparator/U1588  ( .a(\comparator/N459 ), .out(\comparator/n1588 ) );
  inv \comparator/U1587  ( .a(\comparator/N458 ), .out(\comparator/n1587 ) );
  inv \comparator/U1586  ( .a(\comparator/N461 ), .out(\comparator/n1586 ) );
  inv \comparator/U1585  ( .a(\comparator/N460 ), .out(\comparator/n1585 ) );
  inv \comparator/U1584  ( .a(\comparator/N463 ), .out(\comparator/n1584 ) );
  inv \comparator/U1583  ( .a(\comparator/N462 ), .out(\comparator/n1583 ) );
  inv \comparator/U1582  ( .a(\comparator/N465 ), .out(\comparator/n1582 ) );
  inv \comparator/U1581  ( .a(\comparator/N464 ), .out(\comparator/n1581 ) );
  inv \comparator/U1580  ( .a(\comparator/N467 ), .out(\comparator/n1580 ) );
  inv \comparator/U1579  ( .a(\comparator/N466 ), .out(\comparator/n1579 ) );
  inv \comparator/U1578  ( .a(\comparator/N469 ), .out(\comparator/n1578 ) );
  inv \comparator/U1577  ( .a(\comparator/N468 ), .out(\comparator/n1577 ) );
  inv \comparator/U1576  ( .a(\comparator/N471 ), .out(\comparator/n1576 ) );
  inv \comparator/U1575  ( .a(\comparator/N470 ), .out(\comparator/n1575 ) );
  inv \comparator/U1574  ( .a(\comparator/N473 ), .out(\comparator/n1574 ) );
  inv \comparator/U1573  ( .a(\comparator/N472 ), .out(\comparator/n1573 ) );
  inv \comparator/U1572  ( .a(\comparator/N475 ), .out(\comparator/n1572 ) );
  inv \comparator/U1571  ( .a(\comparator/N474 ), .out(\comparator/n1571 ) );
  inv \comparator/U1570  ( .a(\comparator/N477 ), .out(\comparator/n1570 ) );
  inv \comparator/U1569  ( .a(\comparator/N476 ), .out(\comparator/n1569 ) );
  inv \comparator/U1568  ( .a(\comparator/N479 ), .out(\comparator/n1568 ) );
  inv \comparator/U1567  ( .a(\comparator/N478 ), .out(\comparator/n1567 ) );
  inv \comparator/U1566  ( .a(\comparator/N481 ), .out(\comparator/n1566 ) );
  inv \comparator/U1565  ( .a(\comparator/N480 ), .out(\comparator/n1565 ) );
  inv \comparator/U1564  ( .a(\comparator/N483 ), .out(\comparator/n1564 ) );
  inv \comparator/U1563  ( .a(\comparator/N482 ), .out(\comparator/n1563 ) );
  inv \comparator/U1562  ( .a(\comparator/N485 ), .out(\comparator/n1562 ) );
  inv \comparator/U1561  ( .a(\comparator/N484 ), .out(\comparator/n1561 ) );
  inv \comparator/U1560  ( .a(\comparator/N487 ), .out(\comparator/n1560 ) );
  inv \comparator/U1559  ( .a(\comparator/N486 ), .out(\comparator/n1559 ) );
  inv \comparator/U1558  ( .a(\comparator/N489 ), .out(\comparator/n1558 ) );
  inv \comparator/U1557  ( .a(\comparator/N488 ), .out(\comparator/n1557 ) );
  inv \comparator/U1556  ( .a(\comparator/N491 ), .out(\comparator/n1556 ) );
  inv \comparator/U1555  ( .a(\comparator/N490 ), .out(\comparator/n1555 ) );
  inv \comparator/U1554  ( .a(\comparator/N493 ), .out(\comparator/n1554 ) );
  inv \comparator/U1553  ( .a(\comparator/N492 ), .out(\comparator/n1553 ) );
  inv \comparator/U1552  ( .a(\comparator/N495 ), .out(\comparator/n1552 ) );
  inv \comparator/U1551  ( .a(\comparator/N494 ), .out(\comparator/n1551 ) );
  inv \comparator/U1550  ( .a(\comparator/N497 ), .out(\comparator/n1550 ) );
  inv \comparator/U1549  ( .a(\comparator/N496 ), .out(\comparator/n1549 ) );
  inv \comparator/U1548  ( .a(\comparator/N499 ), .out(\comparator/n1548 ) );
  inv \comparator/U1547  ( .a(\comparator/N498 ), .out(\comparator/n1547 ) );
  inv \comparator/U1546  ( .a(\comparator/N501 ), .out(\comparator/n1546 ) );
  inv \comparator/U1545  ( .a(\comparator/N500 ), .out(\comparator/n1545 ) );
  inv \comparator/U1544  ( .a(\comparator/N503 ), .out(\comparator/n1544 ) );
  inv \comparator/U1543  ( .a(\comparator/N502 ), .out(\comparator/n1543 ) );
  inv \comparator/U1542  ( .a(\comparator/N505 ), .out(\comparator/n1542 ) );
  inv \comparator/U1541  ( .a(\comparator/N504 ), .out(\comparator/n1541 ) );
  inv \comparator/U1540  ( .a(\comparator/N507 ), .out(\comparator/n1540 ) );
  inv \comparator/U1539  ( .a(\comparator/N506 ), .out(\comparator/n1539 ) );
  inv \comparator/U1538  ( .a(\comparator/N509 ), .out(\comparator/n1538 ) );
  inv \comparator/U1537  ( .a(\comparator/N508 ), .out(\comparator/n1537 ) );
  inv \comparator/U1536  ( .a(\comparator/N511 ), .out(\comparator/n1536 ) );
  inv \comparator/U1535  ( .a(\comparator/N510 ), .out(\comparator/n1535 ) );
  inv \comparator/U1534  ( .a(\comparator/N513 ), .out(\comparator/n1534 ) );
  inv \comparator/U1533  ( .a(\comparator/N512 ), .out(\comparator/n1533 ) );
  inv \comparator/U1532  ( .a(\comparator/N515 ), .out(\comparator/n1532 ) );
  inv \comparator/U1531  ( .a(\comparator/N514 ), .out(\comparator/n1531 ) );
  inv \comparator/U1530  ( .a(\comparator/N517 ), .out(\comparator/n1530 ) );
  inv \comparator/U1529  ( .a(\comparator/N516 ), .out(\comparator/n1529 ) );
  inv \comparator/U1528  ( .a(\comparator/N519 ), .out(\comparator/n1528 ) );
  inv \comparator/U1527  ( .a(\comparator/N518 ), .out(\comparator/n1527 ) );
  inv \comparator/U1526  ( .a(\comparator/N521 ), .out(\comparator/n1526 ) );
  inv \comparator/U1525  ( .a(\comparator/N520 ), .out(\comparator/n1525 ) );
  inv \comparator/U1524  ( .a(\comparator/N523 ), .out(\comparator/n1524 ) );
  inv \comparator/U1523  ( .a(\comparator/N522 ), .out(\comparator/n1523 ) );
  inv \comparator/U1522  ( .a(\comparator/N525 ), .out(\comparator/n1522 ) );
  inv \comparator/U1521  ( .a(\comparator/N524 ), .out(\comparator/n1521 ) );
  inv \comparator/U1520  ( .a(\comparator/N527 ), .out(\comparator/n1520 ) );
  inv \comparator/U1519  ( .a(\comparator/N526 ), .out(\comparator/n1519 ) );
  inv \comparator/U1518  ( .a(\comparator/N529 ), .out(\comparator/n1518 ) );
  inv \comparator/U1517  ( .a(\comparator/N528 ), .out(\comparator/n1517 ) );
  inv \comparator/U1516  ( .a(\comparator/N531 ), .out(\comparator/n1516 ) );
  inv \comparator/U1515  ( .a(\comparator/N530 ), .out(\comparator/n1515 ) );
  inv \comparator/U1514  ( .a(\comparator/N533 ), .out(\comparator/n1514 ) );
  inv \comparator/U1513  ( .a(\comparator/N532 ), .out(\comparator/n1513 ) );
  inv \comparator/U1512  ( .a(\comparator/N535 ), .out(\comparator/n1512 ) );
  inv \comparator/U1511  ( .a(\comparator/N534 ), .out(\comparator/n1511 ) );
  inv \comparator/U1510  ( .a(\comparator/N537 ), .out(\comparator/n1510 ) );
  inv \comparator/U1509  ( .a(\comparator/N536 ), .out(\comparator/n1509 ) );
  inv \comparator/U1508  ( .a(\comparator/N539 ), .out(\comparator/n1508 ) );
  inv \comparator/U1507  ( .a(\comparator/N538 ), .out(\comparator/n1507 ) );
  inv \comparator/U1506  ( .a(\comparator/N541 ), .out(\comparator/n1506 ) );
  inv \comparator/U1505  ( .a(\comparator/N540 ), .out(\comparator/n1505 ) );
  inv \comparator/U1504  ( .a(\comparator/N543 ), .out(\comparator/n1504 ) );
  inv \comparator/U1503  ( .a(\comparator/N542 ), .out(\comparator/n1503 ) );
  inv \comparator/U1502  ( .a(\comparator/N545 ), .out(\comparator/n1502 ) );
  inv \comparator/U1501  ( .a(\comparator/N544 ), .out(\comparator/n1501 ) );
  inv \comparator/U1500  ( .a(\comparator/N547 ), .out(\comparator/n1500 ) );
  inv \comparator/U1499  ( .a(\comparator/N546 ), .out(\comparator/n1499 ) );
  inv \comparator/U1498  ( .a(\comparator/N549 ), .out(\comparator/n1498 ) );
  inv \comparator/U1497  ( .a(\comparator/N548 ), .out(\comparator/n1497 ) );
  inv \comparator/U1496  ( .a(\comparator/N551 ), .out(\comparator/n1496 ) );
  inv \comparator/U1495  ( .a(\comparator/N550 ), .out(\comparator/n1495 ) );
  inv \comparator/U1494  ( .a(\comparator/N553 ), .out(\comparator/n1494 ) );
  inv \comparator/U1493  ( .a(\comparator/N552 ), .out(\comparator/n1493 ) );
  inv \comparator/U1492  ( .a(\comparator/N555 ), .out(\comparator/n1492 ) );
  inv \comparator/U1491  ( .a(\comparator/N554 ), .out(\comparator/n1491 ) );
  inv \comparator/U1490  ( .a(\comparator/N557 ), .out(\comparator/n1490 ) );
  inv \comparator/U1489  ( .a(\comparator/N556 ), .out(\comparator/n1489 ) );
  inv \comparator/U1488  ( .a(\comparator/N559 ), .out(\comparator/n1488 ) );
  inv \comparator/U1487  ( .a(\comparator/N558 ), .out(\comparator/n1487 ) );
  inv \comparator/U1486  ( .a(\comparator/N561 ), .out(\comparator/n1486 ) );
  inv \comparator/U1485  ( .a(\comparator/N560 ), .out(\comparator/n1485 ) );
  inv \comparator/U1484  ( .a(\comparator/N563 ), .out(\comparator/n1484 ) );
  inv \comparator/U1483  ( .a(\comparator/N562 ), .out(\comparator/n1483 ) );
  inv \comparator/U1482  ( .a(\comparator/N565 ), .out(\comparator/n1482 ) );
  inv \comparator/U1481  ( .a(\comparator/N564 ), .out(\comparator/n1481 ) );
  inv \comparator/U1480  ( .a(\comparator/N567 ), .out(\comparator/n1480 ) );
  inv \comparator/U1479  ( .a(\comparator/N566 ), .out(\comparator/n1479 ) );
  inv \comparator/U1478  ( .a(\comparator/N569 ), .out(\comparator/n1478 ) );
  inv \comparator/U1477  ( .a(\comparator/N568 ), .out(\comparator/n1477 ) );
  inv \comparator/U1476  ( .a(\comparator/N571 ), .out(\comparator/n1476 ) );
  inv \comparator/U1475  ( .a(\comparator/N570 ), .out(\comparator/n1475 ) );
  inv \comparator/U1474  ( .a(\comparator/N573 ), .out(\comparator/n1474 ) );
  inv \comparator/U1473  ( .a(\comparator/N572 ), .out(\comparator/n1473 ) );
  inv \comparator/U1472  ( .a(\comparator/N575 ), .out(\comparator/n1472 ) );
  inv \comparator/U1471  ( .a(\comparator/N574 ), .out(\comparator/n1471 ) );
  inv \comparator/U1470  ( .a(\comparator/N577 ), .out(\comparator/n1470 ) );
  inv \comparator/U1469  ( .a(\comparator/N576 ), .out(\comparator/n1469 ) );
  inv \comparator/U1468  ( .a(\comparator/N579 ), .out(\comparator/n1468 ) );
  inv \comparator/U1467  ( .a(\comparator/N578 ), .out(\comparator/n1467 ) );
  inv \comparator/U1466  ( .a(\comparator/N581 ), .out(\comparator/n1466 ) );
  inv \comparator/U1465  ( .a(\comparator/N580 ), .out(\comparator/n1465 ) );
  inv \comparator/U1464  ( .a(\comparator/N583 ), .out(\comparator/n1464 ) );
  inv \comparator/U1463  ( .a(\comparator/N582 ), .out(\comparator/n1463 ) );
  inv \comparator/U1462  ( .a(\comparator/N585 ), .out(\comparator/n1462 ) );
  inv \comparator/U1461  ( .a(\comparator/N584 ), .out(\comparator/n1461 ) );
  inv \comparator/U1460  ( .a(\comparator/N587 ), .out(\comparator/n1460 ) );
  inv \comparator/U1459  ( .a(\comparator/N586 ), .out(\comparator/n1459 ) );
  inv \comparator/U1458  ( .a(\comparator/N589 ), .out(\comparator/n1458 ) );
  inv \comparator/U1457  ( .a(\comparator/N588 ), .out(\comparator/n1457 ) );
  inv \comparator/U1456  ( .a(\comparator/N591 ), .out(\comparator/n1456 ) );
  inv \comparator/U1455  ( .a(\comparator/N590 ), .out(\comparator/n1455 ) );
  inv \comparator/U1454  ( .a(\comparator/N593 ), .out(\comparator/n1454 ) );
  inv \comparator/U1453  ( .a(\comparator/N592 ), .out(\comparator/n1453 ) );
  inv \comparator/U1452  ( .a(\comparator/N595 ), .out(\comparator/n1452 ) );
  inv \comparator/U1451  ( .a(\comparator/N594 ), .out(\comparator/n1451 ) );
  inv \comparator/U1450  ( .a(\comparator/N597 ), .out(\comparator/n1450 ) );
  inv \comparator/U1449  ( .a(\comparator/N596 ), .out(\comparator/n1449 ) );
  inv \comparator/U1448  ( .a(\comparator/N599 ), .out(\comparator/n1448 ) );
  inv \comparator/U1447  ( .a(\comparator/N598 ), .out(\comparator/n1447 ) );
  inv \comparator/U1446  ( .a(\comparator/N601 ), .out(\comparator/n1446 ) );
  inv \comparator/U1445  ( .a(\comparator/N600 ), .out(\comparator/n1445 ) );
  inv \comparator/U1444  ( .a(\comparator/N603 ), .out(\comparator/n1444 ) );
  inv \comparator/U1443  ( .a(\comparator/N602 ), .out(\comparator/n1443 ) );
  inv \comparator/U1442  ( .a(\comparator/N605 ), .out(\comparator/n1442 ) );
  inv \comparator/U1441  ( .a(\comparator/N604 ), .out(\comparator/n1441 ) );
  inv \comparator/U1440  ( .a(\comparator/N607 ), .out(\comparator/n1440 ) );
  inv \comparator/U1439  ( .a(\comparator/N606 ), .out(\comparator/n1439 ) );
  inv \comparator/U1438  ( .a(\comparator/N609 ), .out(\comparator/n1438 ) );
  inv \comparator/U1437  ( .a(\comparator/N608 ), .out(\comparator/n1437 ) );
  inv \comparator/U1436  ( .a(\comparator/N611 ), .out(\comparator/n1436 ) );
  inv \comparator/U1435  ( .a(\comparator/N610 ), .out(\comparator/n1435 ) );
  inv \comparator/U1434  ( .a(\comparator/N613 ), .out(\comparator/n1434 ) );
  inv \comparator/U1433  ( .a(\comparator/N612 ), .out(\comparator/n1433 ) );
  inv \comparator/U1432  ( .a(\comparator/N615 ), .out(\comparator/n1432 ) );
  inv \comparator/U1431  ( .a(\comparator/N614 ), .out(\comparator/n1431 ) );
  inv \comparator/U1430  ( .a(\comparator/N617 ), .out(\comparator/n1430 ) );
  inv \comparator/U1429  ( .a(\comparator/N616 ), .out(\comparator/n1429 ) );
  inv \comparator/U1428  ( .a(\comparator/N619 ), .out(\comparator/n1428 ) );
  inv \comparator/U1427  ( .a(\comparator/N618 ), .out(\comparator/n1427 ) );
  inv \comparator/U1426  ( .a(\comparator/N621 ), .out(\comparator/n1426 ) );
  inv \comparator/U1425  ( .a(\comparator/N620 ), .out(\comparator/n1425 ) );
  inv \comparator/U1424  ( .a(\comparator/N623 ), .out(\comparator/n1424 ) );
  inv \comparator/U1423  ( .a(\comparator/N622 ), .out(\comparator/n1423 ) );
  inv \comparator/U1422  ( .a(\comparator/N625 ), .out(\comparator/n1422 ) );
  inv \comparator/U1421  ( .a(\comparator/N624 ), .out(\comparator/n1421 ) );
  inv \comparator/U1420  ( .a(\comparator/N627 ), .out(\comparator/n1420 ) );
  inv \comparator/U1419  ( .a(\comparator/N626 ), .out(\comparator/n1419 ) );
  inv \comparator/U1418  ( .a(\comparator/N629 ), .out(\comparator/n1418 ) );
  inv \comparator/U1417  ( .a(\comparator/N628 ), .out(\comparator/n1417 ) );
  inv \comparator/U1416  ( .a(\comparator/N631 ), .out(\comparator/n1416 ) );
  inv \comparator/U1415  ( .a(\comparator/N630 ), .out(\comparator/n1415 ) );
  inv \comparator/U1414  ( .a(\comparator/N633 ), .out(\comparator/n1414 ) );
  inv \comparator/U1413  ( .a(\comparator/N632 ), .out(\comparator/n1413 ) );
  inv \comparator/U1412  ( .a(\comparator/N635 ), .out(\comparator/n1412 ) );
  inv \comparator/U1411  ( .a(\comparator/N634 ), .out(\comparator/n1411 ) );
  inv \comparator/U1410  ( .a(\comparator/N637 ), .out(\comparator/n1410 ) );
  inv \comparator/U1409  ( .a(\comparator/N636 ), .out(\comparator/n1409 ) );
  inv \comparator/U1408  ( .a(\comparator/N639 ), .out(\comparator/n1408 ) );
  inv \comparator/U1407  ( .a(\comparator/N638 ), .out(\comparator/n1407 ) );
  inv \comparator/U1406  ( .a(\comparator/N641 ), .out(\comparator/n1406 ) );
  inv \comparator/U1405  ( .a(\comparator/N640 ), .out(\comparator/n1405 ) );
  inv \comparator/U1404  ( .a(\comparator/N643 ), .out(\comparator/n1404 ) );
  inv \comparator/U1403  ( .a(\comparator/N642 ), .out(\comparator/n1403 ) );
  inv \comparator/U1402  ( .a(\comparator/N645 ), .out(\comparator/n1402 ) );
  inv \comparator/U1401  ( .a(\comparator/N644 ), .out(\comparator/n1401 ) );
  inv \comparator/U1400  ( .a(\comparator/N647 ), .out(\comparator/n1400 ) );
  inv \comparator/U1399  ( .a(\comparator/N646 ), .out(\comparator/n1399 ) );
  inv \comparator/U1398  ( .a(\comparator/N649 ), .out(\comparator/n1398 ) );
  inv \comparator/U1397  ( .a(\comparator/N648 ), .out(\comparator/n1397 ) );
  inv \comparator/U1396  ( .a(\comparator/N651 ), .out(\comparator/n1396 ) );
  inv \comparator/U1395  ( .a(\comparator/N650 ), .out(\comparator/n1395 ) );
  inv \comparator/U1394  ( .a(\comparator/N653 ), .out(\comparator/n1394 ) );
  inv \comparator/U1393  ( .a(\comparator/N652 ), .out(\comparator/n1393 ) );
  inv \comparator/U1392  ( .a(\comparator/N655 ), .out(\comparator/n1392 ) );
  inv \comparator/U1391  ( .a(\comparator/N654 ), .out(\comparator/n1391 ) );
  inv \comparator/U1390  ( .a(\comparator/N657 ), .out(\comparator/n1390 ) );
  inv \comparator/U1389  ( .a(\comparator/N656 ), .out(\comparator/n1389 ) );
  inv \comparator/U1388  ( .a(\comparator/N659 ), .out(\comparator/n1388 ) );
  inv \comparator/U1387  ( .a(\comparator/N658 ), .out(\comparator/n1387 ) );
  inv \comparator/U1386  ( .a(\comparator/N661 ), .out(\comparator/n1386 ) );
  inv \comparator/U1385  ( .a(\comparator/N660 ), .out(\comparator/n1385 ) );
  inv \comparator/U1384  ( .a(\comparator/N663 ), .out(\comparator/n1384 ) );
  inv \comparator/U1383  ( .a(\comparator/N662 ), .out(\comparator/n1383 ) );
  inv \comparator/U1382  ( .a(\comparator/N665 ), .out(\comparator/n1382 ) );
  inv \comparator/U1381  ( .a(\comparator/N664 ), .out(\comparator/n1381 ) );
  inv \comparator/U1380  ( .a(\comparator/N667 ), .out(\comparator/n1380 ) );
  inv \comparator/U1379  ( .a(\comparator/N666 ), .out(\comparator/n1379 ) );
  inv \comparator/U1378  ( .a(\comparator/N669 ), .out(\comparator/n1378 ) );
  inv \comparator/U1377  ( .a(\comparator/N668 ), .out(\comparator/n1377 ) );
  inv \comparator/U1376  ( .a(\comparator/N671 ), .out(\comparator/n1376 ) );
  inv \comparator/U1375  ( .a(\comparator/N670 ), .out(\comparator/n1375 ) );
  inv \comparator/U1374  ( .a(\comparator/N673 ), .out(\comparator/n1374 ) );
  inv \comparator/U1373  ( .a(\comparator/N672 ), .out(\comparator/n1373 ) );
  inv \comparator/U1372  ( .a(\comparator/N675 ), .out(\comparator/n1372 ) );
  inv \comparator/U1371  ( .a(\comparator/N674 ), .out(\comparator/n1371 ) );
  inv \comparator/U1370  ( .a(\comparator/N677 ), .out(\comparator/n1370 ) );
  inv \comparator/U1369  ( .a(\comparator/N676 ), .out(\comparator/n1369 ) );
  inv \comparator/U1368  ( .a(\comparator/N679 ), .out(\comparator/n1368 ) );
  inv \comparator/U1367  ( .a(\comparator/N678 ), .out(\comparator/n1367 ) );
  inv \comparator/U1366  ( .a(\comparator/N681 ), .out(\comparator/n1366 ) );
  inv \comparator/U1365  ( .a(\comparator/N680 ), .out(\comparator/n1365 ) );
  inv \comparator/U1364  ( .a(\comparator/N683 ), .out(\comparator/n1364 ) );
  inv \comparator/U1363  ( .a(\comparator/N682 ), .out(\comparator/n1363 ) );
  inv \comparator/U1362  ( .a(\comparator/N685 ), .out(\comparator/n1362 ) );
  inv \comparator/U1361  ( .a(\comparator/N684 ), .out(\comparator/n1361 ) );
  inv \comparator/U1360  ( .a(\comparator/N687 ), .out(\comparator/n1360 ) );
  inv \comparator/U1359  ( .a(\comparator/N686 ), .out(\comparator/n1359 ) );
  inv \comparator/U1358  ( .a(\comparator/N689 ), .out(\comparator/n1358 ) );
  inv \comparator/U1357  ( .a(\comparator/N688 ), .out(\comparator/n1357 ) );
  inv \comparator/U1356  ( .a(\comparator/N691 ), .out(\comparator/n1356 ) );
  inv \comparator/U1355  ( .a(\comparator/N690 ), .out(\comparator/n1355 ) );
  inv \comparator/U1354  ( .a(\comparator/N693 ), .out(\comparator/n1354 ) );
  inv \comparator/U1353  ( .a(\comparator/N692 ), .out(\comparator/n1353 ) );
  inv \comparator/U1352  ( .a(\comparator/N695 ), .out(\comparator/n1352 ) );
  inv \comparator/U1351  ( .a(\comparator/N694 ), .out(\comparator/n1351 ) );
  inv \comparator/U1350  ( .a(\comparator/N697 ), .out(\comparator/n1350 ) );
  inv \comparator/U1349  ( .a(\comparator/N696 ), .out(\comparator/n1349 ) );
  inv \comparator/U1348  ( .a(\comparator/N699 ), .out(\comparator/n1348 ) );
  inv \comparator/U1347  ( .a(\comparator/N698 ), .out(\comparator/n1347 ) );
  inv \comparator/U1346  ( .a(\comparator/N701 ), .out(\comparator/n1346 ) );
  inv \comparator/U1345  ( .a(\comparator/N700 ), .out(\comparator/n1345 ) );
  inv \comparator/U1344  ( .a(\comparator/N703 ), .out(\comparator/n1344 ) );
  inv \comparator/U1343  ( .a(\comparator/N702 ), .out(\comparator/n1343 ) );
  inv \comparator/U1342  ( .a(\comparator/N705 ), .out(\comparator/n1342 ) );
  inv \comparator/U1341  ( .a(\comparator/N704 ), .out(\comparator/n1341 ) );
  inv \comparator/U1340  ( .a(\comparator/N707 ), .out(\comparator/n1340 ) );
  inv \comparator/U1339  ( .a(\comparator/N706 ), .out(\comparator/n1339 ) );
  inv \comparator/U1338  ( .a(\comparator/N709 ), .out(\comparator/n1338 ) );
  inv \comparator/U1337  ( .a(\comparator/N708 ), .out(\comparator/n1337 ) );
  inv \comparator/U1336  ( .a(\comparator/N711 ), .out(\comparator/n1336 ) );
  inv \comparator/U1335  ( .a(\comparator/N710 ), .out(\comparator/n1335 ) );
  inv \comparator/U1334  ( .a(\comparator/N713 ), .out(\comparator/n1334 ) );
  inv \comparator/U1333  ( .a(\comparator/N712 ), .out(\comparator/n1333 ) );
  inv \comparator/U1332  ( .a(\comparator/N715 ), .out(\comparator/n1332 ) );
  inv \comparator/U1331  ( .a(\comparator/N714 ), .out(\comparator/n1331 ) );
  inv \comparator/U1330  ( .a(\comparator/N717 ), .out(\comparator/n1330 ) );
  inv \comparator/U1329  ( .a(\comparator/N716 ), .out(\comparator/n1329 ) );
  inv \comparator/U1328  ( .a(\comparator/N719 ), .out(\comparator/n1328 ) );
  inv \comparator/U1327  ( .a(\comparator/N718 ), .out(\comparator/n1327 ) );
  inv \comparator/U1326  ( .a(\comparator/N721 ), .out(\comparator/n1326 ) );
  inv \comparator/U1325  ( .a(\comparator/N720 ), .out(\comparator/n1325 ) );
  inv \comparator/U1324  ( .a(\comparator/N723 ), .out(\comparator/n1324 ) );
  inv \comparator/U1323  ( .a(\comparator/N722 ), .out(\comparator/n1323 ) );
  inv \comparator/U1322  ( .a(\comparator/N725 ), .out(\comparator/n1322 ) );
  inv \comparator/U1321  ( .a(\comparator/N724 ), .out(\comparator/n1321 ) );
  inv \comparator/U1320  ( .a(\comparator/N727 ), .out(\comparator/n1320 ) );
  inv \comparator/U1319  ( .a(\comparator/N726 ), .out(\comparator/n1319 ) );
  inv \comparator/U1318  ( .a(\comparator/N729 ), .out(\comparator/n1318 ) );
  inv \comparator/U1317  ( .a(\comparator/N728 ), .out(\comparator/n1317 ) );
  inv \comparator/U1316  ( .a(\comparator/N731 ), .out(\comparator/n1316 ) );
  inv \comparator/U1315  ( .a(\comparator/N730 ), .out(\comparator/n1315 ) );
  inv \comparator/U1314  ( .a(\comparator/N733 ), .out(\comparator/n1314 ) );
  inv \comparator/U1313  ( .a(\comparator/N732 ), .out(\comparator/n1313 ) );
  inv \comparator/U1312  ( .a(\comparator/N735 ), .out(\comparator/n1312 ) );
  inv \comparator/U1311  ( .a(\comparator/N734 ), .out(\comparator/n1311 ) );
  inv \comparator/U1310  ( .a(\comparator/N737 ), .out(\comparator/n1310 ) );
  inv \comparator/U1309  ( .a(\comparator/N736 ), .out(\comparator/n1309 ) );
  inv \comparator/U1308  ( .a(\comparator/N739 ), .out(\comparator/n1308 ) );
  inv \comparator/U1307  ( .a(\comparator/N738 ), .out(\comparator/n1307 ) );
  inv \comparator/U1306  ( .a(\comparator/N741 ), .out(\comparator/n1306 ) );
  inv \comparator/U1305  ( .a(\comparator/N740 ), .out(\comparator/n1305 ) );
  inv \comparator/U1304  ( .a(\comparator/N743 ), .out(\comparator/n1304 ) );
  inv \comparator/U1303  ( .a(\comparator/N742 ), .out(\comparator/n1303 ) );
  inv \comparator/U1302  ( .a(\comparator/N745 ), .out(\comparator/n1302 ) );
  inv \comparator/U1301  ( .a(\comparator/N744 ), .out(\comparator/n1301 ) );
  inv \comparator/U1300  ( .a(\comparator/N747 ), .out(\comparator/n1300 ) );
  inv \comparator/U1299  ( .a(\comparator/N746 ), .out(\comparator/n1299 ) );
  inv \comparator/U1298  ( .a(\comparator/N749 ), .out(\comparator/n1298 ) );
  inv \comparator/U1297  ( .a(\comparator/N748 ), .out(\comparator/n1297 ) );
  inv \comparator/U1296  ( .a(\comparator/N751 ), .out(\comparator/n1296 ) );
  inv \comparator/U1295  ( .a(\comparator/N750 ), .out(\comparator/n1295 ) );
  inv \comparator/U1294  ( .a(\comparator/N753 ), .out(\comparator/n1294 ) );
  inv \comparator/U1293  ( .a(\comparator/N752 ), .out(\comparator/n1293 ) );
  inv \comparator/U1292  ( .a(\comparator/N755 ), .out(\comparator/n1292 ) );
  inv \comparator/U1291  ( .a(\comparator/N754 ), .out(\comparator/n1291 ) );
  inv \comparator/U1290  ( .a(\comparator/N757 ), .out(\comparator/n1290 ) );
  inv \comparator/U1289  ( .a(\comparator/N756 ), .out(\comparator/n1289 ) );
  inv \comparator/U1288  ( .a(\comparator/N759 ), .out(\comparator/n1288 ) );
  inv \comparator/U1287  ( .a(\comparator/N758 ), .out(\comparator/n1287 ) );
  inv \comparator/U1286  ( .a(\comparator/N761 ), .out(\comparator/n1286 ) );
  inv \comparator/U1285  ( .a(\comparator/N760 ), .out(\comparator/n1285 ) );
  inv \comparator/U1284  ( .a(\comparator/N763 ), .out(\comparator/n1284 ) );
  inv \comparator/U1283  ( .a(\comparator/N762 ), .out(\comparator/n1283 ) );
  inv \comparator/U1282  ( .a(\comparator/N765 ), .out(\comparator/n1282 ) );
  inv \comparator/U1281  ( .a(\comparator/N764 ), .out(\comparator/n1281 ) );
  inv \comparator/U1280  ( .a(\comparator/N767 ), .out(\comparator/n1280 ) );
  inv \comparator/U1279  ( .a(\comparator/N766 ), .out(\comparator/n1279 ) );
  inv \comparator/U1278  ( .a(\comparator/N769 ), .out(\comparator/n1278 ) );
  inv \comparator/U1277  ( .a(\comparator/N768 ), .out(\comparator/n1277 ) );
  inv \comparator/U1276  ( .a(\comparator/N771 ), .out(\comparator/n1276 ) );
  inv \comparator/U1275  ( .a(\comparator/N770 ), .out(\comparator/n1275 ) );
  inv \comparator/U1274  ( .a(\comparator/N773 ), .out(\comparator/n1274 ) );
  inv \comparator/U1273  ( .a(\comparator/N772 ), .out(\comparator/n1273 ) );
  inv \comparator/U1272  ( .a(\comparator/N775 ), .out(\comparator/n1272 ) );
  inv \comparator/U1271  ( .a(\comparator/N774 ), .out(\comparator/n1271 ) );
  inv \comparator/U1270  ( .a(\comparator/N777 ), .out(\comparator/n1270 ) );
  inv \comparator/U1269  ( .a(\comparator/N776 ), .out(\comparator/n1269 ) );
  inv \comparator/U1268  ( .a(\comparator/N779 ), .out(\comparator/n1268 ) );
  inv \comparator/U1267  ( .a(\comparator/N778 ), .out(\comparator/n1267 ) );
  inv \comparator/U1266  ( .a(\comparator/N781 ), .out(\comparator/n1266 ) );
  inv \comparator/U1265  ( .a(\comparator/N780 ), .out(\comparator/n1265 ) );
  inv \comparator/U1264  ( .a(\comparator/N783 ), .out(\comparator/n1264 ) );
  inv \comparator/U1263  ( .a(\comparator/N782 ), .out(\comparator/n1263 ) );
  inv \comparator/U1262  ( .a(\comparator/N785 ), .out(\comparator/n1262 ) );
  inv \comparator/U1261  ( .a(\comparator/N784 ), .out(\comparator/n1261 ) );
  inv \comparator/U1260  ( .a(\comparator/N787 ), .out(\comparator/n1260 ) );
  inv \comparator/U1259  ( .a(\comparator/N786 ), .out(\comparator/n1259 ) );
  inv \comparator/U1258  ( .a(\comparator/N789 ), .out(\comparator/n1258 ) );
  inv \comparator/U1257  ( .a(\comparator/N788 ), .out(\comparator/n1257 ) );
  inv \comparator/U1256  ( .a(\comparator/N791 ), .out(\comparator/n1256 ) );
  inv \comparator/U1255  ( .a(\comparator/N790 ), .out(\comparator/n1255 ) );
  inv \comparator/U1254  ( .a(\comparator/N793 ), .out(\comparator/n1254 ) );
  inv \comparator/U1253  ( .a(\comparator/N792 ), .out(\comparator/n1253 ) );
  inv \comparator/U1252  ( .a(\comparator/N795 ), .out(\comparator/n1252 ) );
  inv \comparator/U1251  ( .a(\comparator/N794 ), .out(\comparator/n1251 ) );
  inv \comparator/U1250  ( .a(\comparator/N797 ), .out(\comparator/n1250 ) );
  inv \comparator/U1249  ( .a(\comparator/N796 ), .out(\comparator/n1249 ) );
  inv \comparator/U1248  ( .a(\comparator/N799 ), .out(\comparator/n1248 ) );
  inv \comparator/U1247  ( .a(\comparator/N798 ), .out(\comparator/n1247 ) );
  inv \comparator/U1246  ( .a(\comparator/N801 ), .out(\comparator/n1246 ) );
  inv \comparator/U1245  ( .a(\comparator/N800 ), .out(\comparator/n1245 ) );
  inv \comparator/U1244  ( .a(\comparator/N803 ), .out(\comparator/n1244 ) );
  inv \comparator/U1243  ( .a(\comparator/N802 ), .out(\comparator/n1243 ) );
  inv \comparator/U1242  ( .a(\comparator/N805 ), .out(\comparator/n1242 ) );
  inv \comparator/U1241  ( .a(\comparator/N804 ), .out(\comparator/n1241 ) );
  inv \comparator/U1240  ( .a(\comparator/N807 ), .out(\comparator/n1240 ) );
  inv \comparator/U1239  ( .a(\comparator/N806 ), .out(\comparator/n1239 ) );
  inv \comparator/U1238  ( .a(\comparator/N809 ), .out(\comparator/n1238 ) );
  inv \comparator/U1237  ( .a(\comparator/N808 ), .out(\comparator/n1237 ) );
  inv \comparator/U1236  ( .a(\comparator/N811 ), .out(\comparator/n1236 ) );
  inv \comparator/U1235  ( .a(\comparator/N810 ), .out(\comparator/n1235 ) );
  inv \comparator/U1234  ( .a(\comparator/N813 ), .out(\comparator/n1234 ) );
  inv \comparator/U1233  ( .a(\comparator/N812 ), .out(\comparator/n1233 ) );
  inv \comparator/U1232  ( .a(\comparator/N815 ), .out(\comparator/n1232 ) );
  inv \comparator/U1231  ( .a(\comparator/N814 ), .out(\comparator/n1231 ) );
  inv \comparator/U1230  ( .a(\comparator/N817 ), .out(\comparator/n1230 ) );
  inv \comparator/U1229  ( .a(\comparator/N816 ), .out(\comparator/n1229 ) );
  inv \comparator/U1228  ( .a(\comparator/N819 ), .out(\comparator/n1228 ) );
  inv \comparator/U1227  ( .a(\comparator/N818 ), .out(\comparator/n1227 ) );
  inv \comparator/U1226  ( .a(\comparator/N821 ), .out(\comparator/n1226 ) );
  inv \comparator/U1225  ( .a(\comparator/N820 ), .out(\comparator/n1225 ) );
  inv \comparator/U1224  ( .a(\comparator/N823 ), .out(\comparator/n1224 ) );
  inv \comparator/U1223  ( .a(\comparator/N822 ), .out(\comparator/n1223 ) );
  inv \comparator/U1222  ( .a(\comparator/N825 ), .out(\comparator/n1222 ) );
  inv \comparator/U1221  ( .a(\comparator/N824 ), .out(\comparator/n1221 ) );
  inv \comparator/U1220  ( .a(\comparator/N827 ), .out(\comparator/n1220 ) );
  inv \comparator/U1219  ( .a(\comparator/N826 ), .out(\comparator/n1219 ) );
  inv \comparator/U1218  ( .a(\comparator/N829 ), .out(\comparator/n1218 ) );
  inv \comparator/U1217  ( .a(\comparator/N828 ), .out(\comparator/n1217 ) );
  inv \comparator/U1216  ( .a(\comparator/N831 ), .out(\comparator/n1216 ) );
  inv \comparator/U1215  ( .a(\comparator/N830 ), .out(\comparator/n1215 ) );
  inv \comparator/U1214  ( .a(\comparator/N833 ), .out(\comparator/n1214 ) );
  inv \comparator/U1213  ( .a(\comparator/N832 ), .out(\comparator/n1213 ) );
  inv \comparator/U1212  ( .a(\comparator/N835 ), .out(\comparator/n1212 ) );
  inv \comparator/U1211  ( .a(\comparator/N834 ), .out(\comparator/n1211 ) );
  inv \comparator/U1210  ( .a(\comparator/N837 ), .out(\comparator/n1210 ) );
  inv \comparator/U1209  ( .a(\comparator/N836 ), .out(\comparator/n1209 ) );
  inv \comparator/U1208  ( .a(\comparator/N839 ), .out(\comparator/n1208 ) );
  inv \comparator/U1207  ( .a(\comparator/N838 ), .out(\comparator/n1207 ) );
  inv \comparator/U1206  ( .a(\comparator/N841 ), .out(\comparator/n1206 ) );
  inv \comparator/U1205  ( .a(\comparator/N840 ), .out(\comparator/n1205 ) );
  inv \comparator/U1204  ( .a(\comparator/N843 ), .out(\comparator/n1204 ) );
  inv \comparator/U1203  ( .a(\comparator/N842 ), .out(\comparator/n1203 ) );
  inv \comparator/U1202  ( .a(\comparator/N845 ), .out(\comparator/n1202 ) );
  inv \comparator/U1201  ( .a(\comparator/N844 ), .out(\comparator/n1201 ) );
  inv \comparator/U1200  ( .a(\comparator/N847 ), .out(\comparator/n1200 ) );
  inv \comparator/U1199  ( .a(\comparator/N846 ), .out(\comparator/n1199 ) );
  inv \comparator/U1198  ( .a(\comparator/N849 ), .out(\comparator/n1198 ) );
  inv \comparator/U1197  ( .a(\comparator/N848 ), .out(\comparator/n1197 ) );
  inv \comparator/U1196  ( .a(\comparator/N851 ), .out(\comparator/n1196 ) );
  inv \comparator/U1195  ( .a(\comparator/N850 ), .out(\comparator/n1195 ) );
  inv \comparator/U1194  ( .a(\comparator/N853 ), .out(\comparator/n1194 ) );
  inv \comparator/U1193  ( .a(\comparator/N852 ), .out(\comparator/n1193 ) );
  inv \comparator/U1192  ( .a(\comparator/N855 ), .out(\comparator/n1192 ) );
  inv \comparator/U1191  ( .a(\comparator/N854 ), .out(\comparator/n1191 ) );
  inv \comparator/U1190  ( .a(\comparator/N857 ), .out(\comparator/n1190 ) );
  inv \comparator/U1189  ( .a(\comparator/N856 ), .out(\comparator/n1189 ) );
  inv \comparator/U1188  ( .a(\comparator/N859 ), .out(\comparator/n1188 ) );
  inv \comparator/U1187  ( .a(\comparator/N858 ), .out(\comparator/n1187 ) );
  inv \comparator/U1186  ( .a(\comparator/N861 ), .out(\comparator/n1186 ) );
  inv \comparator/U1185  ( .a(\comparator/N860 ), .out(\comparator/n1185 ) );
  inv \comparator/U1184  ( .a(\comparator/N863 ), .out(\comparator/n1184 ) );
  inv \comparator/U1183  ( .a(\comparator/N862 ), .out(\comparator/n1183 ) );
  inv \comparator/U1182  ( .a(\comparator/N865 ), .out(\comparator/n1182 ) );
  inv \comparator/U1181  ( .a(\comparator/N864 ), .out(\comparator/n1181 ) );
  inv \comparator/U1180  ( .a(\comparator/N867 ), .out(\comparator/n1180 ) );
  inv \comparator/U1179  ( .a(\comparator/N866 ), .out(\comparator/n1179 ) );
  inv \comparator/U1178  ( .a(\comparator/N869 ), .out(\comparator/n1178 ) );
  inv \comparator/U1177  ( .a(\comparator/N868 ), .out(\comparator/n1177 ) );
  inv \comparator/U1176  ( .a(\comparator/N871 ), .out(\comparator/n1176 ) );
  inv \comparator/U1175  ( .a(\comparator/N870 ), .out(\comparator/n1175 ) );
  inv \comparator/U1174  ( .a(\comparator/N873 ), .out(\comparator/n1174 ) );
  inv \comparator/U1173  ( .a(\comparator/N872 ), .out(\comparator/n1173 ) );
  inv \comparator/U1172  ( .a(\comparator/N875 ), .out(\comparator/n1172 ) );
  inv \comparator/U1171  ( .a(\comparator/N874 ), .out(\comparator/n1171 ) );
  inv \comparator/U1170  ( .a(\comparator/N877 ), .out(\comparator/n1170 ) );
  inv \comparator/U1169  ( .a(\comparator/N876 ), .out(\comparator/n1169 ) );
  inv \comparator/U1168  ( .a(\comparator/N879 ), .out(\comparator/n1168 ) );
  inv \comparator/U1167  ( .a(\comparator/N878 ), .out(\comparator/n1167 ) );
  inv \comparator/U1166  ( .a(\comparator/N881 ), .out(\comparator/n1166 ) );
  inv \comparator/U1165  ( .a(\comparator/N880 ), .out(\comparator/n1165 ) );
  inv \comparator/U1164  ( .a(\comparator/N883 ), .out(\comparator/n1164 ) );
  inv \comparator/U1163  ( .a(\comparator/N882 ), .out(\comparator/n1163 ) );
  inv \comparator/U1162  ( .a(\comparator/N885 ), .out(\comparator/n1162 ) );
  inv \comparator/U1161  ( .a(\comparator/N884 ), .out(\comparator/n1161 ) );
  inv \comparator/U1160  ( .a(\comparator/N887 ), .out(\comparator/n1160 ) );
  inv \comparator/U1159  ( .a(\comparator/N886 ), .out(\comparator/n1159 ) );
  inv \comparator/U1158  ( .a(\comparator/N889 ), .out(\comparator/n1158 ) );
  inv \comparator/U1157  ( .a(\comparator/N888 ), .out(\comparator/n1157 ) );
  inv \comparator/U1156  ( .a(\comparator/N891 ), .out(\comparator/n1156 ) );
  inv \comparator/U1155  ( .a(\comparator/N890 ), .out(\comparator/n1155 ) );
  inv \comparator/U1154  ( .a(\comparator/N893 ), .out(\comparator/n1154 ) );
  inv \comparator/U1153  ( .a(\comparator/N892 ), .out(\comparator/n1153 ) );
  inv \comparator/U1152  ( .a(\comparator/N895 ), .out(\comparator/n1152 ) );
  inv \comparator/U1151  ( .a(\comparator/N894 ), .out(\comparator/n1151 ) );
  inv \comparator/U1150  ( .a(\comparator/N897 ), .out(\comparator/n1150 ) );
  inv \comparator/U1149  ( .a(\comparator/N896 ), .out(\comparator/n1149 ) );
  inv \comparator/U1148  ( .a(\comparator/N899 ), .out(\comparator/n1148 ) );
  inv \comparator/U1147  ( .a(\comparator/N898 ), .out(\comparator/n1147 ) );
  inv \comparator/U1146  ( .a(\comparator/N901 ), .out(\comparator/n1146 ) );
  inv \comparator/U1145  ( .a(\comparator/N900 ), .out(\comparator/n1145 ) );
  inv \comparator/U1144  ( .a(\comparator/N903 ), .out(\comparator/n1144 ) );
  inv \comparator/U1143  ( .a(\comparator/N902 ), .out(\comparator/n1143 ) );
  inv \comparator/U1142  ( .a(\comparator/N905 ), .out(\comparator/n1142 ) );
  inv \comparator/U1141  ( .a(\comparator/N904 ), .out(\comparator/n1141 ) );
  inv \comparator/U1140  ( .a(\comparator/N907 ), .out(\comparator/n1140 ) );
  inv \comparator/U1139  ( .a(\comparator/N906 ), .out(\comparator/n1139 ) );
  inv \comparator/U1138  ( .a(\comparator/N909 ), .out(\comparator/n1138 ) );
  inv \comparator/U1137  ( .a(\comparator/N908 ), .out(\comparator/n1137 ) );
  inv \comparator/U1136  ( .a(\comparator/N911 ), .out(\comparator/n1136 ) );
  inv \comparator/U1135  ( .a(\comparator/N910 ), .out(\comparator/n1135 ) );
  inv \comparator/U1134  ( .a(\comparator/N913 ), .out(\comparator/n1134 ) );
  inv \comparator/U1133  ( .a(\comparator/N912 ), .out(\comparator/n1133 ) );
  inv \comparator/U1132  ( .a(\comparator/N915 ), .out(\comparator/n1132 ) );
  inv \comparator/U1131  ( .a(\comparator/N914 ), .out(\comparator/n1131 ) );
  inv \comparator/U1130  ( .a(\comparator/N917 ), .out(\comparator/n1130 ) );
  inv \comparator/U1129  ( .a(\comparator/N916 ), .out(\comparator/n1129 ) );
  inv \comparator/U1128  ( .a(\comparator/N919 ), .out(\comparator/n1128 ) );
  inv \comparator/U1127  ( .a(\comparator/N918 ), .out(\comparator/n1127 ) );
  inv \comparator/U1126  ( .a(\comparator/N921 ), .out(\comparator/n1126 ) );
  inv \comparator/U1125  ( .a(\comparator/N920 ), .out(\comparator/n1125 ) );
  inv \comparator/U1124  ( .a(\comparator/N923 ), .out(\comparator/n1124 ) );
  inv \comparator/U1123  ( .a(\comparator/N922 ), .out(\comparator/n1123 ) );
  inv \comparator/U1122  ( .a(\comparator/N925 ), .out(\comparator/n1122 ) );
  inv \comparator/U1121  ( .a(\comparator/N924 ), .out(\comparator/n1121 ) );
  inv \comparator/U1120  ( .a(\comparator/N927 ), .out(\comparator/n1120 ) );
  inv \comparator/U1119  ( .a(\comparator/N926 ), .out(\comparator/n1119 ) );
  inv \comparator/U1118  ( .a(\comparator/N929 ), .out(\comparator/n1118 ) );
  inv \comparator/U1117  ( .a(\comparator/N928 ), .out(\comparator/n1117 ) );
  inv \comparator/U1116  ( .a(\comparator/N931 ), .out(\comparator/n1116 ) );
  inv \comparator/U1115  ( .a(\comparator/N930 ), .out(\comparator/n1115 ) );
  inv \comparator/U1114  ( .a(\comparator/N933 ), .out(\comparator/n1114 ) );
  inv \comparator/U1113  ( .a(\comparator/N932 ), .out(\comparator/n1113 ) );
  inv \comparator/U1112  ( .a(\comparator/N935 ), .out(\comparator/n1112 ) );
  inv \comparator/U1111  ( .a(\comparator/N934 ), .out(\comparator/n1111 ) );
  inv \comparator/U1110  ( .a(\comparator/N937 ), .out(\comparator/n1110 ) );
  inv \comparator/U1109  ( .a(\comparator/N936 ), .out(\comparator/n1109 ) );
  inv \comparator/U1108  ( .a(\comparator/N939 ), .out(\comparator/n1108 ) );
  inv \comparator/U1107  ( .a(\comparator/N938 ), .out(\comparator/n1107 ) );
  inv \comparator/U1106  ( .a(\comparator/N941 ), .out(\comparator/n1106 ) );
  inv \comparator/U1105  ( .a(\comparator/N940 ), .out(\comparator/n1105 ) );
  inv \comparator/U1104  ( .a(\comparator/N943 ), .out(\comparator/n1104 ) );
  inv \comparator/U1103  ( .a(\comparator/N942 ), .out(\comparator/n1103 ) );
  inv \comparator/U1102  ( .a(\comparator/N945 ), .out(\comparator/n1102 ) );
  inv \comparator/U1101  ( .a(\comparator/N944 ), .out(\comparator/n1101 ) );
  inv \comparator/U1100  ( .a(\comparator/N947 ), .out(\comparator/n1100 ) );
  inv \comparator/U1099  ( .a(\comparator/N946 ), .out(\comparator/n1099 ) );
  inv \comparator/U1098  ( .a(\comparator/N949 ), .out(\comparator/n1098 ) );
  inv \comparator/U1097  ( .a(\comparator/N948 ), .out(\comparator/n1097 ) );
  inv \comparator/U1096  ( .a(\comparator/N951 ), .out(\comparator/n1096 ) );
  inv \comparator/U1095  ( .a(\comparator/N950 ), .out(\comparator/n1095 ) );
  inv \comparator/U1094  ( .a(\comparator/N953 ), .out(\comparator/n1094 ) );
  inv \comparator/U1093  ( .a(\comparator/N952 ), .out(\comparator/n1093 ) );
  inv \comparator/U1092  ( .a(\comparator/N955 ), .out(\comparator/n1092 ) );
  inv \comparator/U1091  ( .a(\comparator/N954 ), .out(\comparator/n1091 ) );
  inv \comparator/U1090  ( .a(\comparator/N957 ), .out(\comparator/n1090 ) );
  inv \comparator/U1089  ( .a(\comparator/N956 ), .out(\comparator/n1089 ) );
  inv \comparator/U1088  ( .a(\comparator/N959 ), .out(\comparator/n1088 ) );
  inv \comparator/U1087  ( .a(\comparator/N958 ), .out(\comparator/n1087 ) );
  inv \comparator/U1086  ( .a(\comparator/N961 ), .out(\comparator/n1086 ) );
  inv \comparator/U1085  ( .a(\comparator/N960 ), .out(\comparator/n1085 ) );
  inv \comparator/U1084  ( .a(\comparator/N963 ), .out(\comparator/n1084 ) );
  inv \comparator/U1083  ( .a(\comparator/N962 ), .out(\comparator/n1083 ) );
  inv \comparator/U1082  ( .a(\comparator/N965 ), .out(\comparator/n1082 ) );
  inv \comparator/U1081  ( .a(\comparator/N964 ), .out(\comparator/n1081 ) );
  inv \comparator/U1080  ( .a(\comparator/N967 ), .out(\comparator/n1080 ) );
  inv \comparator/U1079  ( .a(\comparator/N966 ), .out(\comparator/n1079 ) );
  inv \comparator/U1078  ( .a(\comparator/N969 ), .out(\comparator/n1078 ) );
  inv \comparator/U1077  ( .a(\comparator/N968 ), .out(\comparator/n1077 ) );
  inv \comparator/U1076  ( .a(\comparator/N971 ), .out(\comparator/n1076 ) );
  inv \comparator/U1075  ( .a(\comparator/N970 ), .out(\comparator/n1075 ) );
  inv \comparator/U1074  ( .a(\comparator/N973 ), .out(\comparator/n1074 ) );
  inv \comparator/U1073  ( .a(\comparator/N972 ), .out(\comparator/n1073 ) );
  inv \comparator/U1072  ( .a(\comparator/N975 ), .out(\comparator/n1072 ) );
  inv \comparator/U1071  ( .a(\comparator/N974 ), .out(\comparator/n1071 ) );
  inv \comparator/U1070  ( .a(\comparator/N977 ), .out(\comparator/n1070 ) );
  inv \comparator/U1069  ( .a(\comparator/N976 ), .out(\comparator/n1069 ) );
  inv \comparator/U1068  ( .a(\comparator/N979 ), .out(\comparator/n1068 ) );
  inv \comparator/U1067  ( .a(\comparator/N978 ), .out(\comparator/n1067 ) );
  inv \comparator/U1066  ( .a(\comparator/N981 ), .out(\comparator/n1066 ) );
  inv \comparator/U1065  ( .a(\comparator/N980 ), .out(\comparator/n1065 ) );
  inv \comparator/U1064  ( .a(\comparator/N983 ), .out(\comparator/n1064 ) );
  inv \comparator/U1063  ( .a(\comparator/N982 ), .out(\comparator/n1063 ) );
  inv \comparator/U1062  ( .a(\comparator/N985 ), .out(\comparator/n1062 ) );
  inv \comparator/U1061  ( .a(\comparator/N984 ), .out(\comparator/n1061 ) );
  inv \comparator/U1060  ( .a(\comparator/N987 ), .out(\comparator/n1060 ) );
  inv \comparator/U1059  ( .a(\comparator/N986 ), .out(\comparator/n1059 ) );
  inv \comparator/U1058  ( .a(\comparator/N989 ), .out(\comparator/n1058 ) );
  inv \comparator/U1057  ( .a(\comparator/N988 ), .out(\comparator/n1057 ) );
  inv \comparator/U1056  ( .a(\comparator/N991 ), .out(\comparator/n1056 ) );
  inv \comparator/U1055  ( .a(\comparator/N990 ), .out(\comparator/n1055 ) );
  inv \comparator/U1054  ( .a(\comparator/N993 ), .out(\comparator/n1054 ) );
  inv \comparator/U1053  ( .a(\comparator/N992 ), .out(\comparator/n1053 ) );
  inv \comparator/U1052  ( .a(\comparator/N995 ), .out(\comparator/n1052 ) );
  inv \comparator/U1051  ( .a(\comparator/N994 ), .out(\comparator/n1051 ) );
  inv \comparator/U1050  ( .a(\comparator/N997 ), .out(\comparator/n1050 ) );
  inv \comparator/U1049  ( .a(\comparator/N996 ), .out(\comparator/n1049 ) );
  inv \comparator/U1048  ( .a(\comparator/N999 ), .out(\comparator/n1048 ) );
  inv \comparator/U1047  ( .a(\comparator/N998 ), .out(\comparator/n1047 ) );
  inv \comparator/U1046  ( .a(\comparator/N1001 ), .out(\comparator/n1046 )
         );
  inv \comparator/U1045  ( .a(\comparator/N1000 ), .out(\comparator/n1045 )
         );
  inv \comparator/U1044  ( .a(\comparator/N1003 ), .out(\comparator/n1044 )
         );
  inv \comparator/U1043  ( .a(\comparator/N1002 ), .out(\comparator/n1043 )
         );
  inv \comparator/U1042  ( .a(\comparator/N1005 ), .out(\comparator/n1042 )
         );
  inv \comparator/U1041  ( .a(\comparator/N1004 ), .out(\comparator/n1041 )
         );
  inv \comparator/U1040  ( .a(\comparator/N1007 ), .out(\comparator/n1040 )
         );
  inv \comparator/U1039  ( .a(\comparator/N1006 ), .out(\comparator/n1039 )
         );
  inv \comparator/U1038  ( .a(\comparator/N1009 ), .out(\comparator/n1038 )
         );
  inv \comparator/U1037  ( .a(\comparator/N1008 ), .out(\comparator/n1037 )
         );
  inv \comparator/U1036  ( .a(\comparator/N1011 ), .out(\comparator/n1036 )
         );
  inv \comparator/U1035  ( .a(\comparator/N1010 ), .out(\comparator/n1035 )
         );
  inv \comparator/U1034  ( .a(\comparator/N1013 ), .out(\comparator/n1034 )
         );
  inv \comparator/U1033  ( .a(\comparator/N1012 ), .out(\comparator/n1033 )
         );
  inv \comparator/U1032  ( .a(\comparator/N1015 ), .out(\comparator/n1032 )
         );
  inv \comparator/U1031  ( .a(\comparator/N1014 ), .out(\comparator/n1031 )
         );
  inv \comparator/U1030  ( .a(\comparator/N1017 ), .out(\comparator/n1030 )
         );
  inv \comparator/U1029  ( .a(\comparator/N1016 ), .out(\comparator/n1029 )
         );
  inv \comparator/U1028  ( .a(\comparator/N1019 ), .out(\comparator/n1028 )
         );
  inv \comparator/U1027  ( .a(\comparator/N1018 ), .out(\comparator/n1027 )
         );
  inv \comparator/U1026  ( .a(\comparator/N1021 ), .out(\comparator/n1026 )
         );
  inv \comparator/U1025  ( .a(\comparator/N1020 ), .out(\comparator/n1025 )
         );
  inv \comparator/U1024  ( .a(\comparator/N1023 ), .out(\comparator/n1024 )
         );
  inv \comparator/U1023  ( .a(\comparator/N1022 ), .out(\comparator/n1023 )
         );
  inv \comparator/U1022  ( .a(\comparator/N1025 ), .out(\comparator/n1022 )
         );
  inv \comparator/U1021  ( .a(\comparator/N1024 ), .out(\comparator/n1021 )
         );
  inv \comparator/U1020  ( .a(\comparator/N1027 ), .out(\comparator/n1020 )
         );
  inv \comparator/U1019  ( .a(\comparator/N1026 ), .out(\comparator/n1019 )
         );
  inv \comparator/U1018  ( .a(\comparator/N1029 ), .out(\comparator/n1018 )
         );
  inv \comparator/U1017  ( .a(\comparator/N1028 ), .out(\comparator/n1017 )
         );
  inv \comparator/U1016  ( .a(\comparator/N1031 ), .out(\comparator/n1016 )
         );
  inv \comparator/U1015  ( .a(\comparator/N1030 ), .out(\comparator/n1015 )
         );
  inv \comparator/U1014  ( .a(\comparator/N1033 ), .out(\comparator/n1014 )
         );
  inv \comparator/U1013  ( .a(\comparator/N1032 ), .out(\comparator/n1013 )
         );
  inv \comparator/U1012  ( .a(\comparator/N1035 ), .out(\comparator/n1012 )
         );
  inv \comparator/U1011  ( .a(\comparator/N1034 ), .out(\comparator/n1011 )
         );
  inv \comparator/U1010  ( .a(\comparator/N1037 ), .out(\comparator/n1010 )
         );
  inv \comparator/U1009  ( .a(\comparator/N1036 ), .out(\comparator/n1009 )
         );
  inv \comparator/U1008  ( .a(\comparator/N1039 ), .out(\comparator/n1008 )
         );
  inv \comparator/U1007  ( .a(\comparator/N1038 ), .out(\comparator/n1007 )
         );
  inv \comparator/U1006  ( .a(\comparator/N1041 ), .out(\comparator/n1006 )
         );
  inv \comparator/U1005  ( .a(\comparator/N1040 ), .out(\comparator/n1005 )
         );
  inv \comparator/U1004  ( .a(\comparator/N1043 ), .out(\comparator/n1004 )
         );
  inv \comparator/U1003  ( .a(\comparator/N1042 ), .out(\comparator/n1003 )
         );
  inv \comparator/U1002  ( .a(\comparator/N1045 ), .out(\comparator/n1002 )
         );
  inv \comparator/U1001  ( .a(\comparator/N1044 ), .out(\comparator/n1001 )
         );
  inv \comparator/U1000  ( .a(\comparator/N1047 ), .out(\comparator/n1000 )
         );
  inv \comparator/U999  ( .a(\comparator/N1046 ), .out(\comparator/n999 ) );
  inv \comparator/U998  ( .a(\comparator/N1049 ), .out(\comparator/n998 ) );
  inv \comparator/U997  ( .a(\comparator/N1048 ), .out(\comparator/n997 ) );
  inv \comparator/U996  ( .a(\comparator/N1051 ), .out(\comparator/n996 ) );
  inv \comparator/U995  ( .a(\comparator/N1050 ), .out(\comparator/n995 ) );
  inv \comparator/U994  ( .a(\comparator/N1053 ), .out(\comparator/n994 ) );
  inv \comparator/U993  ( .a(\comparator/N1052 ), .out(\comparator/n993 ) );
  inv \comparator/U992  ( .a(\comparator/N1055 ), .out(\comparator/n992 ) );
  inv \comparator/U991  ( .a(\comparator/N1054 ), .out(\comparator/n991 ) );
  inv \comparator/U990  ( .a(\comparator/N1057 ), .out(\comparator/n990 ) );
  inv \comparator/U989  ( .a(\comparator/N1056 ), .out(\comparator/n989 ) );
  inv \comparator/U988  ( .a(\comparator/N1059 ), .out(\comparator/n988 ) );
  inv \comparator/U987  ( .a(\comparator/N1058 ), .out(\comparator/n987 ) );
  inv \comparator/U986  ( .a(\comparator/N1061 ), .out(\comparator/n986 ) );
  inv \comparator/U985  ( .a(\comparator/N1060 ), .out(\comparator/n985 ) );
  inv \comparator/U984  ( .a(\comparator/N1063 ), .out(\comparator/n984 ) );
  inv \comparator/U983  ( .a(\comparator/N1062 ), .out(\comparator/n983 ) );
  inv \comparator/U982  ( .a(\comparator/N1065 ), .out(\comparator/n982 ) );
  inv \comparator/U981  ( .a(\comparator/N1064 ), .out(\comparator/n981 ) );
  inv \comparator/U980  ( .a(\comparator/N1067 ), .out(\comparator/n980 ) );
  inv \comparator/U979  ( .a(\comparator/N1066 ), .out(\comparator/n979 ) );
  inv \comparator/U978  ( .a(\comparator/N1069 ), .out(\comparator/n978 ) );
  inv \comparator/U977  ( .a(\comparator/N1068 ), .out(\comparator/n977 ) );
  inv \comparator/U976  ( .a(\comparator/N1071 ), .out(\comparator/n976 ) );
  inv \comparator/U975  ( .a(\comparator/N1070 ), .out(\comparator/n975 ) );
  inv \comparator/U974  ( .a(\comparator/N1073 ), .out(\comparator/n974 ) );
  inv \comparator/U973  ( .a(\comparator/N1072 ), .out(\comparator/n973 ) );
  inv \comparator/U972  ( .a(\comparator/N1075 ), .out(\comparator/n972 ) );
  inv \comparator/U971  ( .a(\comparator/N1074 ), .out(\comparator/n971 ) );
  inv \comparator/U970  ( .a(\comparator/N1077 ), .out(\comparator/n970 ) );
  inv \comparator/U969  ( .a(\comparator/N1076 ), .out(\comparator/n969 ) );
  inv \comparator/U968  ( .a(\comparator/N1079 ), .out(\comparator/n968 ) );
  inv \comparator/U967  ( .a(\comparator/N1078 ), .out(\comparator/n967 ) );
  inv \comparator/U966  ( .a(\comparator/N1081 ), .out(\comparator/n966 ) );
  inv \comparator/U965  ( .a(\comparator/N1080 ), .out(\comparator/n965 ) );
  inv \comparator/U964  ( .a(\comparator/N1083 ), .out(\comparator/n964 ) );
  inv \comparator/U963  ( .a(\comparator/N1082 ), .out(\comparator/n963 ) );
  inv \comparator/U962  ( .a(\comparator/N1085 ), .out(\comparator/n962 ) );
  inv \comparator/U961  ( .a(\comparator/N1084 ), .out(\comparator/n961 ) );
  inv \comparator/U960  ( .a(\comparator/N1087 ), .out(\comparator/n960 ) );
  inv \comparator/U959  ( .a(\comparator/N1086 ), .out(\comparator/n959 ) );
  inv \comparator/U958  ( .a(\comparator/N1089 ), .out(\comparator/n958 ) );
  inv \comparator/U957  ( .a(\comparator/N1088 ), .out(\comparator/n957 ) );
  inv \comparator/U956  ( .a(\comparator/N1091 ), .out(\comparator/n956 ) );
  inv \comparator/U955  ( .a(\comparator/N1090 ), .out(\comparator/n955 ) );
  inv \comparator/U954  ( .a(\comparator/N1093 ), .out(\comparator/n954 ) );
  inv \comparator/U953  ( .a(\comparator/N1092 ), .out(\comparator/n953 ) );
  inv \comparator/U952  ( .a(\comparator/N1095 ), .out(\comparator/n952 ) );
  inv \comparator/U951  ( .a(\comparator/N1094 ), .out(\comparator/n951 ) );
  inv \comparator/U950  ( .a(\comparator/N1097 ), .out(\comparator/n950 ) );
  inv \comparator/U949  ( .a(\comparator/N1096 ), .out(\comparator/n949 ) );
  inv \comparator/U948  ( .a(\comparator/N1099 ), .out(\comparator/n948 ) );
  inv \comparator/U947  ( .a(\comparator/N1098 ), .out(\comparator/n947 ) );
  inv \comparator/U946  ( .a(\comparator/N1101 ), .out(\comparator/n946 ) );
  inv \comparator/U945  ( .a(\comparator/N1100 ), .out(\comparator/n945 ) );
  inv \comparator/U944  ( .a(\comparator/N1103 ), .out(\comparator/n944 ) );
  inv \comparator/U943  ( .a(\comparator/N1102 ), .out(\comparator/n943 ) );
  inv \comparator/U942  ( .a(\comparator/N1105 ), .out(\comparator/n942 ) );
  inv \comparator/U941  ( .a(\comparator/N1104 ), .out(\comparator/n941 ) );
  inv \comparator/U940  ( .a(\comparator/N1107 ), .out(\comparator/n940 ) );
  inv \comparator/U939  ( .a(\comparator/N1106 ), .out(\comparator/n939 ) );
  inv \comparator/U938  ( .a(\comparator/N1109 ), .out(\comparator/n938 ) );
  inv \comparator/U937  ( .a(\comparator/N1108 ), .out(\comparator/n937 ) );
  inv \comparator/U936  ( .a(\comparator/N1111 ), .out(\comparator/n936 ) );
  inv \comparator/U935  ( .a(\comparator/N1110 ), .out(\comparator/n935 ) );
  inv \comparator/U934  ( .a(\comparator/N1113 ), .out(\comparator/n934 ) );
  inv \comparator/U933  ( .a(\comparator/N1112 ), .out(\comparator/n933 ) );
  inv \comparator/U932  ( .a(\comparator/N1115 ), .out(\comparator/n932 ) );
  inv \comparator/U931  ( .a(\comparator/N1114 ), .out(\comparator/n931 ) );
  inv \comparator/U930  ( .a(\comparator/N1117 ), .out(\comparator/n930 ) );
  inv \comparator/U929  ( .a(\comparator/N1116 ), .out(\comparator/n929 ) );
  inv \comparator/U928  ( .a(\comparator/N1119 ), .out(\comparator/n928 ) );
  inv \comparator/U927  ( .a(\comparator/N1118 ), .out(\comparator/n927 ) );
  inv \comparator/U926  ( .a(\comparator/N1121 ), .out(\comparator/n926 ) );
  inv \comparator/U925  ( .a(\comparator/N1120 ), .out(\comparator/n925 ) );
  inv \comparator/U924  ( .a(\comparator/N1123 ), .out(\comparator/n924 ) );
  inv \comparator/U923  ( .a(\comparator/N1122 ), .out(\comparator/n923 ) );
  inv \comparator/U922  ( .a(\comparator/N1125 ), .out(\comparator/n922 ) );
  inv \comparator/U921  ( .a(\comparator/N1124 ), .out(\comparator/n921 ) );
  inv \comparator/U920  ( .a(\comparator/N1127 ), .out(\comparator/n920 ) );
  inv \comparator/U919  ( .a(\comparator/N1126 ), .out(\comparator/n919 ) );
  inv \comparator/U918  ( .a(\comparator/N1129 ), .out(\comparator/n918 ) );
  inv \comparator/U917  ( .a(\comparator/N1128 ), .out(\comparator/n917 ) );
  inv \comparator/U916  ( .a(\comparator/N1131 ), .out(\comparator/n916 ) );
  inv \comparator/U915  ( .a(\comparator/N1130 ), .out(\comparator/n915 ) );
  inv \comparator/U914  ( .a(\comparator/N1133 ), .out(\comparator/n914 ) );
  inv \comparator/U913  ( .a(\comparator/N1132 ), .out(\comparator/n913 ) );
  inv \comparator/U912  ( .a(\comparator/N1135 ), .out(\comparator/n912 ) );
  inv \comparator/U911  ( .a(\comparator/N1134 ), .out(\comparator/n911 ) );
  inv \comparator/U910  ( .a(\comparator/N1137 ), .out(\comparator/n910 ) );
  inv \comparator/U909  ( .a(\comparator/N1136 ), .out(\comparator/n909 ) );
  inv \comparator/U908  ( .a(\comparator/N1139 ), .out(\comparator/n908 ) );
  inv \comparator/U907  ( .a(\comparator/N1138 ), .out(\comparator/n907 ) );
  inv \comparator/U906  ( .a(\comparator/N1141 ), .out(\comparator/n906 ) );
  inv \comparator/U905  ( .a(\comparator/N1140 ), .out(\comparator/n905 ) );
  inv \comparator/U904  ( .a(\comparator/N1143 ), .out(\comparator/n904 ) );
  inv \comparator/U903  ( .a(\comparator/N1142 ), .out(\comparator/n903 ) );
  inv \comparator/U902  ( .a(\comparator/N1145 ), .out(\comparator/n902 ) );
  inv \comparator/U901  ( .a(\comparator/N1144 ), .out(\comparator/n901 ) );
  inv \comparator/U900  ( .a(\comparator/N1147 ), .out(\comparator/n900 ) );
  inv \comparator/U899  ( .a(\comparator/N1146 ), .out(\comparator/n899 ) );
  inv \comparator/U898  ( .a(\comparator/N1149 ), .out(\comparator/n898 ) );
  inv \comparator/U897  ( .a(\comparator/N1148 ), .out(\comparator/n897 ) );
  inv \comparator/U896  ( .a(\comparator/N1151 ), .out(\comparator/n896 ) );
  inv \comparator/U895  ( .a(\comparator/N1150 ), .out(\comparator/n895 ) );
  inv \comparator/U894  ( .a(\comparator/N1153 ), .out(\comparator/n894 ) );
  inv \comparator/U893  ( .a(\comparator/N1152 ), .out(\comparator/n893 ) );
  inv \comparator/U892  ( .a(\comparator/N1155 ), .out(\comparator/n892 ) );
  inv \comparator/U891  ( .a(\comparator/N1154 ), .out(\comparator/n891 ) );
  inv \comparator/U890  ( .a(\comparator/N1157 ), .out(\comparator/n890 ) );
  inv \comparator/U889  ( .a(\comparator/N1156 ), .out(\comparator/n889 ) );
  inv \comparator/U888  ( .a(\comparator/N1159 ), .out(\comparator/n888 ) );
  inv \comparator/U887  ( .a(\comparator/N1158 ), .out(\comparator/n887 ) );
  inv \comparator/U886  ( .a(\comparator/N1161 ), .out(\comparator/n886 ) );
  inv \comparator/U885  ( .a(\comparator/N1160 ), .out(\comparator/n885 ) );
  inv \comparator/U884  ( .a(\comparator/N1163 ), .out(\comparator/n884 ) );
  inv \comparator/U883  ( .a(\comparator/N1162 ), .out(\comparator/n883 ) );
  inv \comparator/U882  ( .a(\comparator/N1165 ), .out(\comparator/n882 ) );
  inv \comparator/U881  ( .a(\comparator/N1164 ), .out(\comparator/n881 ) );
  inv \comparator/U880  ( .a(\comparator/N1167 ), .out(\comparator/n880 ) );
  inv \comparator/U879  ( .a(\comparator/N1166 ), .out(\comparator/n879 ) );
  inv \comparator/U878  ( .a(\comparator/N1169 ), .out(\comparator/n878 ) );
  inv \comparator/U877  ( .a(\comparator/N1168 ), .out(\comparator/n877 ) );
  inv \comparator/U876  ( .a(\comparator/N1171 ), .out(\comparator/n876 ) );
  inv \comparator/U875  ( .a(\comparator/N1170 ), .out(\comparator/n875 ) );
  inv \comparator/U874  ( .a(\comparator/N1173 ), .out(\comparator/n874 ) );
  inv \comparator/U873  ( .a(\comparator/N1172 ), .out(\comparator/n873 ) );
  inv \comparator/U872  ( .a(\comparator/N1175 ), .out(\comparator/n872 ) );
  inv \comparator/U871  ( .a(\comparator/N1174 ), .out(\comparator/n871 ) );
  inv \comparator/U870  ( .a(\comparator/N1177 ), .out(\comparator/n870 ) );
  inv \comparator/U869  ( .a(\comparator/N1176 ), .out(\comparator/n869 ) );
  inv \comparator/U868  ( .a(\comparator/N1179 ), .out(\comparator/n868 ) );
  inv \comparator/U867  ( .a(\comparator/N1178 ), .out(\comparator/n867 ) );
  inv \comparator/U866  ( .a(\comparator/N1181 ), .out(\comparator/n866 ) );
  inv \comparator/U865  ( .a(\comparator/N1180 ), .out(\comparator/n865 ) );
  inv \comparator/U864  ( .a(\comparator/N1183 ), .out(\comparator/n864 ) );
  inv \comparator/U863  ( .a(\comparator/N1182 ), .out(\comparator/n863 ) );
  inv \comparator/U862  ( .a(\comparator/N1185 ), .out(\comparator/n862 ) );
  inv \comparator/U861  ( .a(\comparator/N1184 ), .out(\comparator/n861 ) );
  inv \comparator/U860  ( .a(\comparator/N1187 ), .out(\comparator/n860 ) );
  inv \comparator/U859  ( .a(\comparator/N1186 ), .out(\comparator/n859 ) );
  inv \comparator/U858  ( .a(\comparator/N1189 ), .out(\comparator/n858 ) );
  inv \comparator/U857  ( .a(\comparator/N1188 ), .out(\comparator/n857 ) );
  inv \comparator/U856  ( .a(\comparator/N1191 ), .out(\comparator/n856 ) );
  inv \comparator/U855  ( .a(\comparator/N1190 ), .out(\comparator/n855 ) );
  inv \comparator/U854  ( .a(\comparator/N1193 ), .out(\comparator/n854 ) );
  inv \comparator/U853  ( .a(\comparator/N1192 ), .out(\comparator/n853 ) );
  inv \comparator/U852  ( .a(\comparator/N1195 ), .out(\comparator/n852 ) );
  inv \comparator/U851  ( .a(\comparator/N1194 ), .out(\comparator/n851 ) );
  inv \comparator/U850  ( .a(\comparator/N1197 ), .out(\comparator/n850 ) );
  inv \comparator/U849  ( .a(\comparator/N1196 ), .out(\comparator/n849 ) );
  inv \comparator/U848  ( .a(\comparator/N1199 ), .out(\comparator/n848 ) );
  inv \comparator/U847  ( .a(\comparator/N1198 ), .out(\comparator/n847 ) );
  inv \comparator/U846  ( .a(\comparator/N1201 ), .out(\comparator/n846 ) );
  inv \comparator/U845  ( .a(\comparator/N1200 ), .out(\comparator/n845 ) );
  inv \comparator/U844  ( .a(\comparator/N1203 ), .out(\comparator/n844 ) );
  inv \comparator/U843  ( .a(\comparator/N1202 ), .out(\comparator/n843 ) );
  inv \comparator/U842  ( .a(\comparator/N1205 ), .out(\comparator/n842 ) );
  inv \comparator/U841  ( .a(\comparator/N1204 ), .out(\comparator/n841 ) );
  inv \comparator/U840  ( .a(\comparator/N1207 ), .out(\comparator/n840 ) );
  inv \comparator/U839  ( .a(\comparator/N1206 ), .out(\comparator/n839 ) );
  inv \comparator/U838  ( .a(\comparator/N1209 ), .out(\comparator/n838 ) );
  inv \comparator/U837  ( .a(\comparator/N1208 ), .out(\comparator/n837 ) );
  inv \comparator/U836  ( .a(\comparator/N1211 ), .out(\comparator/n836 ) );
  inv \comparator/U835  ( .a(\comparator/N1210 ), .out(\comparator/n835 ) );
  inv \comparator/U834  ( .a(\comparator/N1213 ), .out(\comparator/n834 ) );
  inv \comparator/U833  ( .a(\comparator/N1212 ), .out(\comparator/n833 ) );
  inv \comparator/U832  ( .a(\comparator/N1215 ), .out(\comparator/n832 ) );
  inv \comparator/U831  ( .a(\comparator/N1214 ), .out(\comparator/n831 ) );
  inv \comparator/U830  ( .a(\comparator/N1217 ), .out(\comparator/n830 ) );
  inv \comparator/U829  ( .a(\comparator/N1216 ), .out(\comparator/n829 ) );
  inv \comparator/U828  ( .a(\comparator/N1219 ), .out(\comparator/n828 ) );
  inv \comparator/U827  ( .a(\comparator/N1218 ), .out(\comparator/n827 ) );
  inv \comparator/U826  ( .a(\comparator/N1221 ), .out(\comparator/n826 ) );
  inv \comparator/U825  ( .a(\comparator/N1220 ), .out(\comparator/n825 ) );
  inv \comparator/U824  ( .a(\comparator/N1223 ), .out(\comparator/n824 ) );
  inv \comparator/U823  ( .a(\comparator/N1222 ), .out(\comparator/n823 ) );
  inv \comparator/U822  ( .a(\comparator/N1225 ), .out(\comparator/n822 ) );
  inv \comparator/U821  ( .a(\comparator/N1224 ), .out(\comparator/n821 ) );
  inv \comparator/U820  ( .a(\comparator/N1227 ), .out(\comparator/n820 ) );
  inv \comparator/U819  ( .a(\comparator/N1226 ), .out(\comparator/n819 ) );
  inv \comparator/U818  ( .a(\comparator/N1229 ), .out(\comparator/n818 ) );
  inv \comparator/U817  ( .a(\comparator/N1228 ), .out(\comparator/n817 ) );
  inv \comparator/U816  ( .a(\comparator/N1231 ), .out(\comparator/n816 ) );
  inv \comparator/U815  ( .a(\comparator/N1230 ), .out(\comparator/n815 ) );
  inv \comparator/U814  ( .a(\comparator/N1233 ), .out(\comparator/n814 ) );
  inv \comparator/U813  ( .a(\comparator/N1232 ), .out(\comparator/n813 ) );
  inv \comparator/U812  ( .a(\comparator/N1235 ), .out(\comparator/n812 ) );
  inv \comparator/U811  ( .a(\comparator/N1234 ), .out(\comparator/n811 ) );
  inv \comparator/U810  ( .a(\comparator/N1237 ), .out(\comparator/n810 ) );
  inv \comparator/U809  ( .a(\comparator/N1236 ), .out(\comparator/n809 ) );
  inv \comparator/U808  ( .a(\comparator/N1239 ), .out(\comparator/n808 ) );
  inv \comparator/U807  ( .a(\comparator/N1238 ), .out(\comparator/n807 ) );
  inv \comparator/U806  ( .a(\comparator/N1241 ), .out(\comparator/n806 ) );
  inv \comparator/U805  ( .a(\comparator/N1240 ), .out(\comparator/n805 ) );
  inv \comparator/U804  ( .a(\comparator/N1243 ), .out(\comparator/n804 ) );
  inv \comparator/U803  ( .a(\comparator/N1242 ), .out(\comparator/n803 ) );
  inv \comparator/U802  ( .a(\comparator/N1245 ), .out(\comparator/n802 ) );
  inv \comparator/U801  ( .a(\comparator/N1244 ), .out(\comparator/n801 ) );
  inv \comparator/U800  ( .a(\comparator/N1247 ), .out(\comparator/n800 ) );
  inv \comparator/U799  ( .a(\comparator/N1246 ), .out(\comparator/n799 ) );
  inv \comparator/U798  ( .a(\comparator/N1249 ), .out(\comparator/n798 ) );
  inv \comparator/U797  ( .a(\comparator/N1248 ), .out(\comparator/n797 ) );
  inv \comparator/U796  ( .a(\comparator/N1251 ), .out(\comparator/n796 ) );
  inv \comparator/U795  ( .a(\comparator/N1250 ), .out(\comparator/n795 ) );
  inv \comparator/U794  ( .a(\comparator/N1253 ), .out(\comparator/n794 ) );
  inv \comparator/U793  ( .a(\comparator/N1252 ), .out(\comparator/n793 ) );
  inv \comparator/U792  ( .a(\comparator/N1255 ), .out(\comparator/n792 ) );
  inv \comparator/U791  ( .a(\comparator/N1254 ), .out(\comparator/n791 ) );
  inv \comparator/U790  ( .a(\comparator/N1257 ), .out(\comparator/n790 ) );
  inv \comparator/U789  ( .a(\comparator/N1256 ), .out(\comparator/n789 ) );
  inv \comparator/U788  ( .a(\comparator/N1259 ), .out(\comparator/n788 ) );
  inv \comparator/U787  ( .a(\comparator/N1258 ), .out(\comparator/n787 ) );
  inv \comparator/U786  ( .a(\comparator/N1261 ), .out(\comparator/n786 ) );
  inv \comparator/U785  ( .a(\comparator/N1260 ), .out(\comparator/n785 ) );
  inv \comparator/U784  ( .a(\comparator/N1263 ), .out(\comparator/n784 ) );
  inv \comparator/U783  ( .a(\comparator/N1262 ), .out(\comparator/n783 ) );
  inv \comparator/U782  ( .a(\comparator/N1265 ), .out(\comparator/n782 ) );
  inv \comparator/U781  ( .a(\comparator/N1264 ), .out(\comparator/n781 ) );
  inv \comparator/U780  ( .a(\comparator/N1267 ), .out(\comparator/n780 ) );
  inv \comparator/U779  ( .a(\comparator/N1266 ), .out(\comparator/n779 ) );
  inv \comparator/U778  ( .a(\comparator/N1269 ), .out(\comparator/n778 ) );
  inv \comparator/U777  ( .a(\comparator/N1268 ), .out(\comparator/n777 ) );
  inv \comparator/U776  ( .a(\comparator/N1271 ), .out(\comparator/n776 ) );
  inv \comparator/U775  ( .a(\comparator/N1270 ), .out(\comparator/n775 ) );
  inv \comparator/U774  ( .a(\comparator/N1273 ), .out(\comparator/n774 ) );
  inv \comparator/U773  ( .a(\comparator/N1272 ), .out(\comparator/n773 ) );
  inv \comparator/U772  ( .a(\comparator/N1275 ), .out(\comparator/n772 ) );
  inv \comparator/U771  ( .a(\comparator/N1274 ), .out(\comparator/n771 ) );
  inv \comparator/U770  ( .a(\comparator/N1277 ), .out(\comparator/n770 ) );
  inv \comparator/U769  ( .a(\comparator/N1276 ), .out(\comparator/n769 ) );
  inv \comparator/U768  ( .a(\comparator/N1279 ), .out(\comparator/n768 ) );
  inv \comparator/U767  ( .a(\comparator/N1278 ), .out(\comparator/n767 ) );
  inv \comparator/U766  ( .a(\comparator/N1281 ), .out(\comparator/n766 ) );
  inv \comparator/U765  ( .a(\comparator/N1280 ), .out(\comparator/n765 ) );
  inv \comparator/U764  ( .a(\comparator/N1283 ), .out(\comparator/n764 ) );
  inv \comparator/U763  ( .a(\comparator/N1282 ), .out(\comparator/n763 ) );
  inv \comparator/U762  ( .a(\comparator/N1285 ), .out(\comparator/n762 ) );
  inv \comparator/U761  ( .a(\comparator/N1284 ), .out(\comparator/n761 ) );
  inv \comparator/U760  ( .a(\comparator/N1287 ), .out(\comparator/n760 ) );
  inv \comparator/U759  ( .a(\comparator/N1286 ), .out(\comparator/n759 ) );
  inv \comparator/U758  ( .a(\comparator/N1289 ), .out(\comparator/n758 ) );
  inv \comparator/U757  ( .a(\comparator/N1288 ), .out(\comparator/n757 ) );
  inv \comparator/U756  ( .a(\comparator/N1291 ), .out(\comparator/n756 ) );
  inv \comparator/U755  ( .a(\comparator/N1290 ), .out(\comparator/n755 ) );
  inv \comparator/U754  ( .a(\comparator/N1293 ), .out(\comparator/n754 ) );
  inv \comparator/U753  ( .a(\comparator/N1292 ), .out(\comparator/n753 ) );
  inv \comparator/U752  ( .a(\comparator/N1295 ), .out(\comparator/n752 ) );
  inv \comparator/U751  ( .a(\comparator/N1294 ), .out(\comparator/n751 ) );
  inv \comparator/U750  ( .a(\comparator/N1297 ), .out(\comparator/n750 ) );
  inv \comparator/U749  ( .a(\comparator/N1296 ), .out(\comparator/n749 ) );
  inv \comparator/U748  ( .a(\comparator/N1299 ), .out(\comparator/n748 ) );
  inv \comparator/U747  ( .a(\comparator/N1298 ), .out(\comparator/n747 ) );
  inv \comparator/U746  ( .a(\comparator/N1301 ), .out(\comparator/n746 ) );
  inv \comparator/U745  ( .a(\comparator/N1300 ), .out(\comparator/n745 ) );
  inv \comparator/U744  ( .a(\comparator/N1303 ), .out(\comparator/n744 ) );
  inv \comparator/U743  ( .a(\comparator/N1302 ), .out(\comparator/n743 ) );
  inv \comparator/U742  ( .a(\comparator/N1305 ), .out(\comparator/n742 ) );
  inv \comparator/U741  ( .a(\comparator/N1304 ), .out(\comparator/n741 ) );
  inv \comparator/U740  ( .a(\comparator/N1307 ), .out(\comparator/n740 ) );
  inv \comparator/U739  ( .a(\comparator/N1306 ), .out(\comparator/n739 ) );
  inv \comparator/U738  ( .a(\comparator/N1309 ), .out(\comparator/n738 ) );
  inv \comparator/U737  ( .a(\comparator/N1308 ), .out(\comparator/n737 ) );
  inv \comparator/U736  ( .a(\comparator/N1311 ), .out(\comparator/n736 ) );
  inv \comparator/U735  ( .a(\comparator/N1310 ), .out(\comparator/n735 ) );
  inv \comparator/U734  ( .a(\comparator/N1313 ), .out(\comparator/n734 ) );
  inv \comparator/U733  ( .a(\comparator/N1312 ), .out(\comparator/n733 ) );
  inv \comparator/U732  ( .a(\comparator/N1315 ), .out(\comparator/n732 ) );
  inv \comparator/U731  ( .a(\comparator/N1314 ), .out(\comparator/n731 ) );
  inv \comparator/U730  ( .a(\comparator/N1317 ), .out(\comparator/n730 ) );
  inv \comparator/U729  ( .a(\comparator/N1316 ), .out(\comparator/n729 ) );
  inv \comparator/U728  ( .a(\comparator/N1319 ), .out(\comparator/n728 ) );
  inv \comparator/U727  ( .a(\comparator/N1318 ), .out(\comparator/n727 ) );
  inv \comparator/U726  ( .a(\comparator/N1321 ), .out(\comparator/n726 ) );
  inv \comparator/U725  ( .a(\comparator/N1320 ), .out(\comparator/n725 ) );
  inv \comparator/U724  ( .a(\comparator/N1323 ), .out(\comparator/n724 ) );
  inv \comparator/U723  ( .a(\comparator/N1322 ), .out(\comparator/n723 ) );
  inv \comparator/U722  ( .a(\comparator/N1325 ), .out(\comparator/n722 ) );
  inv \comparator/U721  ( .a(\comparator/N1324 ), .out(\comparator/n721 ) );
  inv \comparator/U720  ( .a(\comparator/N1327 ), .out(\comparator/n720 ) );
  inv \comparator/U719  ( .a(\comparator/N1326 ), .out(\comparator/n719 ) );
  inv \comparator/U718  ( .a(\comparator/N1329 ), .out(\comparator/n718 ) );
  inv \comparator/U717  ( .a(\comparator/N1328 ), .out(\comparator/n717 ) );
  inv \comparator/U716  ( .a(\comparator/N1331 ), .out(\comparator/n716 ) );
  inv \comparator/U715  ( .a(\comparator/N1330 ), .out(\comparator/n715 ) );
  inv \comparator/U714  ( .a(\comparator/N1333 ), .out(\comparator/n714 ) );
  inv \comparator/U713  ( .a(\comparator/N1332 ), .out(\comparator/n713 ) );
  inv \comparator/U712  ( .a(\comparator/N1335 ), .out(\comparator/n712 ) );
  inv \comparator/U711  ( .a(\comparator/N1334 ), .out(\comparator/n711 ) );
  inv \comparator/U710  ( .a(\comparator/N1337 ), .out(\comparator/n710 ) );
  inv \comparator/U709  ( .a(\comparator/N1336 ), .out(\comparator/n709 ) );
  inv \comparator/U708  ( .a(\comparator/N1339 ), .out(\comparator/n708 ) );
  inv \comparator/U707  ( .a(\comparator/N1338 ), .out(\comparator/n707 ) );
  inv \comparator/U706  ( .a(\comparator/N1341 ), .out(\comparator/n706 ) );
  inv \comparator/U705  ( .a(\comparator/N1340 ), .out(\comparator/n705 ) );
  inv \comparator/U704  ( .a(\comparator/N1343 ), .out(\comparator/n704 ) );
  inv \comparator/U703  ( .a(\comparator/N1342 ), .out(\comparator/n703 ) );
  inv \comparator/U702  ( .a(\comparator/N1345 ), .out(\comparator/n702 ) );
  inv \comparator/U701  ( .a(\comparator/N1344 ), .out(\comparator/n701 ) );
  inv \comparator/U700  ( .a(\comparator/N1347 ), .out(\comparator/n700 ) );
  inv \comparator/U699  ( .a(\comparator/N1346 ), .out(\comparator/n699 ) );
  inv \comparator/U698  ( .a(\comparator/N1349 ), .out(\comparator/n698 ) );
  inv \comparator/U697  ( .a(\comparator/N1348 ), .out(\comparator/n697 ) );
  inv \comparator/U696  ( .a(\comparator/N1351 ), .out(\comparator/n696 ) );
  inv \comparator/U695  ( .a(\comparator/N1350 ), .out(\comparator/n695 ) );
  inv \comparator/U694  ( .a(\comparator/N1353 ), .out(\comparator/n694 ) );
  inv \comparator/U693  ( .a(\comparator/N1352 ), .out(\comparator/n693 ) );
  inv \comparator/U692  ( .a(\comparator/N1355 ), .out(\comparator/n692 ) );
  inv \comparator/U691  ( .a(\comparator/N1354 ), .out(\comparator/n691 ) );
  inv \comparator/U690  ( .a(\comparator/N1357 ), .out(\comparator/n690 ) );
  inv \comparator/U689  ( .a(\comparator/N1356 ), .out(\comparator/n689 ) );
  inv \comparator/U688  ( .a(\comparator/N1359 ), .out(\comparator/n688 ) );
  inv \comparator/U687  ( .a(\comparator/N1358 ), .out(\comparator/n687 ) );
  inv \comparator/U686  ( .a(\comparator/N1361 ), .out(\comparator/n686 ) );
  inv \comparator/U685  ( .a(\comparator/N1360 ), .out(\comparator/n685 ) );
  inv \comparator/U684  ( .a(\comparator/N1363 ), .out(\comparator/n684 ) );
  inv \comparator/U683  ( .a(\comparator/N1362 ), .out(\comparator/n683 ) );
  inv \comparator/U682  ( .a(\comparator/N1365 ), .out(\comparator/n682 ) );
  inv \comparator/U681  ( .a(\comparator/N1364 ), .out(\comparator/n681 ) );
  inv \comparator/U680  ( .a(\comparator/N1367 ), .out(\comparator/n680 ) );
  inv \comparator/U679  ( .a(\comparator/N1366 ), .out(\comparator/n679 ) );
  inv \comparator/U678  ( .a(\comparator/N1369 ), .out(\comparator/n678 ) );
  inv \comparator/U677  ( .a(\comparator/N1368 ), .out(\comparator/n677 ) );
  inv \comparator/U676  ( .a(\comparator/N1371 ), .out(\comparator/n676 ) );
  inv \comparator/U675  ( .a(\comparator/N1370 ), .out(\comparator/n675 ) );
  inv \comparator/U674  ( .a(\comparator/N1373 ), .out(\comparator/n674 ) );
  inv \comparator/U673  ( .a(\comparator/N1372 ), .out(\comparator/n673 ) );
  inv \comparator/U672  ( .a(\comparator/N1375 ), .out(\comparator/n672 ) );
  inv \comparator/U671  ( .a(\comparator/N1374 ), .out(\comparator/n671 ) );
  inv \comparator/U670  ( .a(\comparator/N1377 ), .out(\comparator/n670 ) );
  inv \comparator/U669  ( .a(\comparator/N1376 ), .out(\comparator/n669 ) );
  inv \comparator/U668  ( .a(\comparator/N1379 ), .out(\comparator/n668 ) );
  inv \comparator/U667  ( .a(\comparator/N1378 ), .out(\comparator/n667 ) );
  inv \comparator/U666  ( .a(\comparator/N1381 ), .out(\comparator/n666 ) );
  inv \comparator/U665  ( .a(\comparator/N1380 ), .out(\comparator/n665 ) );
  inv \comparator/U664  ( .a(\comparator/N1383 ), .out(\comparator/n664 ) );
  inv \comparator/U663  ( .a(\comparator/N1382 ), .out(\comparator/n663 ) );
  inv \comparator/U662  ( .a(\comparator/N1385 ), .out(\comparator/n662 ) );
  inv \comparator/U661  ( .a(\comparator/N1384 ), .out(\comparator/n661 ) );
  inv \comparator/U660  ( .a(\comparator/N1387 ), .out(\comparator/n660 ) );
  inv \comparator/U659  ( .a(\comparator/N1386 ), .out(\comparator/n659 ) );
  inv \comparator/U658  ( .a(\comparator/N1389 ), .out(\comparator/n658 ) );
  inv \comparator/U657  ( .a(\comparator/N1388 ), .out(\comparator/n657 ) );
  inv \comparator/U656  ( .a(\comparator/N1391 ), .out(\comparator/n656 ) );
  inv \comparator/U655  ( .a(\comparator/N1390 ), .out(\comparator/n655 ) );
  inv \comparator/U654  ( .a(\comparator/N1393 ), .out(\comparator/n654 ) );
  inv \comparator/U653  ( .a(\comparator/N1392 ), .out(\comparator/n653 ) );
  inv \comparator/U652  ( .a(\comparator/N1395 ), .out(\comparator/n652 ) );
  inv \comparator/U651  ( .a(\comparator/N1394 ), .out(\comparator/n651 ) );
  inv \comparator/U650  ( .a(\comparator/N1397 ), .out(\comparator/n650 ) );
  inv \comparator/U649  ( .a(\comparator/N1396 ), .out(\comparator/n649 ) );
  inv \comparator/U648  ( .a(\comparator/N1399 ), .out(\comparator/n648 ) );
  inv \comparator/U647  ( .a(\comparator/N1398 ), .out(\comparator/n647 ) );
  inv \comparator/U646  ( .a(\comparator/N1401 ), .out(\comparator/n646 ) );
  inv \comparator/U645  ( .a(\comparator/N1400 ), .out(\comparator/n645 ) );
  inv \comparator/U644  ( .a(\comparator/N1403 ), .out(\comparator/n644 ) );
  inv \comparator/U643  ( .a(\comparator/N1402 ), .out(\comparator/n643 ) );
  inv \comparator/U642  ( .a(\comparator/N1405 ), .out(\comparator/n642 ) );
  inv \comparator/U641  ( .a(\comparator/N1404 ), .out(\comparator/n641 ) );
  inv \comparator/U640  ( .a(\comparator/N1407 ), .out(\comparator/n640 ) );
  inv \comparator/U639  ( .a(\comparator/N1406 ), .out(\comparator/n639 ) );
  inv \comparator/U638  ( .a(\comparator/N1409 ), .out(\comparator/n638 ) );
  inv \comparator/U637  ( .a(\comparator/N1408 ), .out(\comparator/n637 ) );
  inv \comparator/U636  ( .a(\comparator/N1411 ), .out(\comparator/n636 ) );
  inv \comparator/U635  ( .a(\comparator/N1410 ), .out(\comparator/n635 ) );
  inv \comparator/U634  ( .a(\comparator/N1413 ), .out(\comparator/n634 ) );
  inv \comparator/U633  ( .a(\comparator/N1412 ), .out(\comparator/n633 ) );
  inv \comparator/U632  ( .a(\comparator/N1415 ), .out(\comparator/n632 ) );
  inv \comparator/U631  ( .a(\comparator/N1414 ), .out(\comparator/n631 ) );
  inv \comparator/U630  ( .a(\comparator/N1417 ), .out(\comparator/n630 ) );
  inv \comparator/U629  ( .a(\comparator/N1416 ), .out(\comparator/n629 ) );
  inv \comparator/U628  ( .a(\comparator/N1419 ), .out(\comparator/n628 ) );
  inv \comparator/U627  ( .a(\comparator/N1418 ), .out(\comparator/n627 ) );
  inv \comparator/U626  ( .a(\comparator/N1421 ), .out(\comparator/n626 ) );
  inv \comparator/U625  ( .a(\comparator/N1420 ), .out(\comparator/n625 ) );
  inv \comparator/U624  ( .a(\comparator/N1423 ), .out(\comparator/n624 ) );
  inv \comparator/U623  ( .a(\comparator/N1422 ), .out(\comparator/n623 ) );
  inv \comparator/U622  ( .a(\comparator/N1425 ), .out(\comparator/n622 ) );
  inv \comparator/U621  ( .a(\comparator/N1424 ), .out(\comparator/n621 ) );
  inv \comparator/U620  ( .a(\comparator/N1427 ), .out(\comparator/n620 ) );
  inv \comparator/U619  ( .a(\comparator/N1426 ), .out(\comparator/n619 ) );
  inv \comparator/U618  ( .a(\comparator/N1429 ), .out(\comparator/n618 ) );
  inv \comparator/U617  ( .a(\comparator/N1428 ), .out(\comparator/n617 ) );
  inv \comparator/U616  ( .a(\comparator/N1431 ), .out(\comparator/n616 ) );
  inv \comparator/U615  ( .a(\comparator/N1430 ), .out(\comparator/n615 ) );
  inv \comparator/U614  ( .a(\comparator/N1433 ), .out(\comparator/n614 ) );
  inv \comparator/U613  ( .a(\comparator/N1432 ), .out(\comparator/n613 ) );
  inv \comparator/U612  ( .a(\comparator/N1435 ), .out(\comparator/n612 ) );
  inv \comparator/U611  ( .a(\comparator/N1434 ), .out(\comparator/n611 ) );
  inv \comparator/U610  ( .a(\comparator/N1437 ), .out(\comparator/n610 ) );
  inv \comparator/U609  ( .a(\comparator/N1436 ), .out(\comparator/n609 ) );
  inv \comparator/U608  ( .a(\comparator/N1439 ), .out(\comparator/n608 ) );
  inv \comparator/U607  ( .a(\comparator/N1438 ), .out(\comparator/n607 ) );
  inv \comparator/U606  ( .a(\comparator/N1441 ), .out(\comparator/n606 ) );
  inv \comparator/U605  ( .a(\comparator/N1440 ), .out(\comparator/n605 ) );
  inv \comparator/U604  ( .a(\comparator/N1443 ), .out(\comparator/n604 ) );
  inv \comparator/U603  ( .a(\comparator/N1442 ), .out(\comparator/n603 ) );
  inv \comparator/U602  ( .a(\comparator/N1445 ), .out(\comparator/n602 ) );
  inv \comparator/U601  ( .a(\comparator/N1444 ), .out(\comparator/n601 ) );
  inv \comparator/U600  ( .a(\comparator/N1447 ), .out(\comparator/n600 ) );
  inv \comparator/U599  ( .a(\comparator/N1446 ), .out(\comparator/n599 ) );
  inv \comparator/U598  ( .a(\comparator/N1449 ), .out(\comparator/n598 ) );
  inv \comparator/U597  ( .a(\comparator/N1448 ), .out(\comparator/n597 ) );
  inv \comparator/U596  ( .a(\comparator/N1451 ), .out(\comparator/n596 ) );
  inv \comparator/U595  ( .a(\comparator/N1450 ), .out(\comparator/n595 ) );
  inv \comparator/U594  ( .a(\comparator/N1453 ), .out(\comparator/n594 ) );
  inv \comparator/U593  ( .a(\comparator/N1452 ), .out(\comparator/n593 ) );
  inv \comparator/U592  ( .a(\comparator/N1455 ), .out(\comparator/n592 ) );
  inv \comparator/U591  ( .a(\comparator/N1454 ), .out(\comparator/n591 ) );
  inv \comparator/U590  ( .a(\comparator/N1457 ), .out(\comparator/n590 ) );
  inv \comparator/U589  ( .a(\comparator/N1456 ), .out(\comparator/n589 ) );
  inv \comparator/U588  ( .a(\comparator/N1459 ), .out(\comparator/n588 ) );
  inv \comparator/U587  ( .a(\comparator/N1458 ), .out(\comparator/n587 ) );
  inv \comparator/U586  ( .a(\comparator/N1461 ), .out(\comparator/n586 ) );
  inv \comparator/U585  ( .a(\comparator/N1460 ), .out(\comparator/n585 ) );
  inv \comparator/U584  ( .a(\comparator/N1463 ), .out(\comparator/n584 ) );
  inv \comparator/U583  ( .a(\comparator/N1462 ), .out(\comparator/n583 ) );
  inv \comparator/U582  ( .a(\comparator/N1465 ), .out(\comparator/n582 ) );
  inv \comparator/U581  ( .a(\comparator/N1464 ), .out(\comparator/n581 ) );
  inv \comparator/U580  ( .a(\comparator/N1467 ), .out(\comparator/n580 ) );
  inv \comparator/U579  ( .a(\comparator/N1466 ), .out(\comparator/n579 ) );
  inv \comparator/U578  ( .a(\comparator/N1469 ), .out(\comparator/n578 ) );
  inv \comparator/U577  ( .a(\comparator/N1468 ), .out(\comparator/n577 ) );
  inv \comparator/U576  ( .a(\comparator/N1471 ), .out(\comparator/n576 ) );
  inv \comparator/U575  ( .a(\comparator/N1470 ), .out(\comparator/n575 ) );
  inv \comparator/U574  ( .a(\comparator/N1473 ), .out(\comparator/n574 ) );
  inv \comparator/U573  ( .a(\comparator/N1472 ), .out(\comparator/n573 ) );
  inv \comparator/U572  ( .a(\comparator/N1475 ), .out(\comparator/n572 ) );
  inv \comparator/U571  ( .a(\comparator/N1474 ), .out(\comparator/n571 ) );
  inv \comparator/U570  ( .a(\comparator/N1477 ), .out(\comparator/n570 ) );
  inv \comparator/U569  ( .a(\comparator/N1476 ), .out(\comparator/n569 ) );
  inv \comparator/U568  ( .a(\comparator/N1479 ), .out(\comparator/n568 ) );
  inv \comparator/U567  ( .a(\comparator/N1478 ), .out(\comparator/n567 ) );
  inv \comparator/U566  ( .a(\comparator/N1481 ), .out(\comparator/n566 ) );
  inv \comparator/U565  ( .a(\comparator/N1480 ), .out(\comparator/n565 ) );
  inv \comparator/U564  ( .a(\comparator/N1483 ), .out(\comparator/n564 ) );
  inv \comparator/U563  ( .a(\comparator/N1482 ), .out(\comparator/n563 ) );
  inv \comparator/U562  ( .a(\comparator/N1485 ), .out(\comparator/n562 ) );
  inv \comparator/U561  ( .a(\comparator/N1484 ), .out(\comparator/n561 ) );
  inv \comparator/U560  ( .a(\comparator/N1487 ), .out(\comparator/n560 ) );
  inv \comparator/U559  ( .a(\comparator/N1486 ), .out(\comparator/n559 ) );
  inv \comparator/U558  ( .a(\comparator/N1489 ), .out(\comparator/n558 ) );
  inv \comparator/U557  ( .a(\comparator/N1488 ), .out(\comparator/n557 ) );
  inv \comparator/U556  ( .a(\comparator/N1491 ), .out(\comparator/n556 ) );
  inv \comparator/U555  ( .a(\comparator/N1490 ), .out(\comparator/n555 ) );
  inv \comparator/U554  ( .a(\comparator/N1493 ), .out(\comparator/n554 ) );
  inv \comparator/U553  ( .a(\comparator/N1492 ), .out(\comparator/n553 ) );
  inv \comparator/U552  ( .a(\comparator/N1495 ), .out(\comparator/n552 ) );
  inv \comparator/U551  ( .a(\comparator/N1494 ), .out(\comparator/n551 ) );
  inv \comparator/U550  ( .a(\comparator/N1497 ), .out(\comparator/n550 ) );
  inv \comparator/U549  ( .a(\comparator/N1496 ), .out(\comparator/n549 ) );
  inv \comparator/U548  ( .a(\comparator/N1499 ), .out(\comparator/n548 ) );
  inv \comparator/U547  ( .a(\comparator/N1498 ), .out(\comparator/n547 ) );
  inv \comparator/U546  ( .a(\comparator/N1501 ), .out(\comparator/n546 ) );
  inv \comparator/U545  ( .a(\comparator/N1500 ), .out(\comparator/n545 ) );
  inv \comparator/U544  ( .a(\comparator/N1503 ), .out(\comparator/n544 ) );
  inv \comparator/U543  ( .a(\comparator/N1502 ), .out(\comparator/n543 ) );
  inv \comparator/U542  ( .a(\comparator/N1505 ), .out(\comparator/n542 ) );
  inv \comparator/U541  ( .a(\comparator/N1504 ), .out(\comparator/n541 ) );
  inv \comparator/U540  ( .a(\comparator/N1507 ), .out(\comparator/n540 ) );
  inv \comparator/U539  ( .a(\comparator/N1506 ), .out(\comparator/n539 ) );
  inv \comparator/U538  ( .a(\comparator/N1509 ), .out(\comparator/n538 ) );
  inv \comparator/U537  ( .a(\comparator/N1508 ), .out(\comparator/n537 ) );
  inv \comparator/U536  ( .a(\comparator/N1511 ), .out(\comparator/n536 ) );
  inv \comparator/U535  ( .a(\comparator/N1510 ), .out(\comparator/n535 ) );
  inv \comparator/U534  ( .a(\comparator/N1513 ), .out(\comparator/n534 ) );
  inv \comparator/U533  ( .a(\comparator/N1512 ), .out(\comparator/n533 ) );
  inv \comparator/U532  ( .a(\comparator/N1515 ), .out(\comparator/n532 ) );
  inv \comparator/U531  ( .a(\comparator/N1514 ), .out(\comparator/n531 ) );
  inv \comparator/U530  ( .a(\comparator/N1517 ), .out(\comparator/n530 ) );
  inv \comparator/U529  ( .a(\comparator/N1516 ), .out(\comparator/n529 ) );
  inv \comparator/U528  ( .a(\comparator/N1519 ), .out(\comparator/n528 ) );
  inv \comparator/U527  ( .a(\comparator/N1518 ), .out(\comparator/n527 ) );
  inv \comparator/U526  ( .a(\comparator/N1521 ), .out(\comparator/n526 ) );
  inv \comparator/U525  ( .a(\comparator/N1520 ), .out(\comparator/n525 ) );
  inv \comparator/U524  ( .a(\comparator/N1523 ), .out(\comparator/n524 ) );
  inv \comparator/U523  ( .a(\comparator/N1522 ), .out(\comparator/n523 ) );
  inv \comparator/U522  ( .a(\comparator/N1525 ), .out(\comparator/n522 ) );
  inv \comparator/U521  ( .a(\comparator/N1524 ), .out(\comparator/n521 ) );
  inv \comparator/U520  ( .a(\comparator/N1527 ), .out(\comparator/n520 ) );
  inv \comparator/U519  ( .a(\comparator/N1526 ), .out(\comparator/n519 ) );
  inv \comparator/U518  ( .a(\comparator/N1529 ), .out(\comparator/n518 ) );
  inv \comparator/U517  ( .a(\comparator/N1528 ), .out(\comparator/n517 ) );
  inv \comparator/U516  ( .a(\comparator/N1531 ), .out(\comparator/n516 ) );
  inv \comparator/U515  ( .a(\comparator/N1530 ), .out(\comparator/n515 ) );
  inv \comparator/U514  ( .a(\comparator/N1533 ), .out(\comparator/n514 ) );
  inv \comparator/U513  ( .a(\comparator/N1532 ), .out(\comparator/n513 ) );
  inv \comparator/U512  ( .a(\comparator/N1535 ), .out(\comparator/n512 ) );
  inv \comparator/U511  ( .a(\comparator/N1534 ), .out(\comparator/n511 ) );
  inv \comparator/U510  ( .a(\comparator/N1537 ), .out(\comparator/n510 ) );
  inv \comparator/U509  ( .a(\comparator/N1536 ), .out(\comparator/n509 ) );
  inv \comparator/U508  ( .a(\comparator/N1539 ), .out(\comparator/n508 ) );
  inv \comparator/U507  ( .a(\comparator/N1538 ), .out(\comparator/n507 ) );
  inv \comparator/U506  ( .a(\comparator/N1541 ), .out(\comparator/n506 ) );
  inv \comparator/U505  ( .a(\comparator/N1540 ), .out(\comparator/n505 ) );
  inv \comparator/U504  ( .a(\comparator/N1543 ), .out(\comparator/n504 ) );
  inv \comparator/U503  ( .a(\comparator/N1542 ), .out(\comparator/n503 ) );
  inv \comparator/U502  ( .a(\comparator/N1545 ), .out(\comparator/n502 ) );
  inv \comparator/U501  ( .a(\comparator/N1544 ), .out(\comparator/n501 ) );
  inv \comparator/U500  ( .a(\comparator/N1547 ), .out(\comparator/n500 ) );
  inv \comparator/U499  ( .a(\comparator/N1546 ), .out(\comparator/n499 ) );
  inv \comparator/U498  ( .a(\comparator/N1549 ), .out(\comparator/n498 ) );
  inv \comparator/U497  ( .a(\comparator/N1548 ), .out(\comparator/n497 ) );
  inv \comparator/U496  ( .a(\comparator/N1551 ), .out(\comparator/n496 ) );
  inv \comparator/U495  ( .a(\comparator/N1550 ), .out(\comparator/n495 ) );
  inv \comparator/U494  ( .a(\comparator/N1553 ), .out(\comparator/n494 ) );
  inv \comparator/U493  ( .a(\comparator/N1552 ), .out(\comparator/n493 ) );
  inv \comparator/U492  ( .a(\comparator/N1555 ), .out(\comparator/n492 ) );
  inv \comparator/U491  ( .a(\comparator/N1554 ), .out(\comparator/n491 ) );
  inv \comparator/U490  ( .a(\comparator/N1557 ), .out(\comparator/n490 ) );
  inv \comparator/U489  ( .a(\comparator/N1556 ), .out(\comparator/n489 ) );
  inv \comparator/U488  ( .a(\comparator/N1559 ), .out(\comparator/n488 ) );
  inv \comparator/U487  ( .a(\comparator/N1558 ), .out(\comparator/n487 ) );
  inv \comparator/U486  ( .a(\comparator/N1561 ), .out(\comparator/n486 ) );
  inv \comparator/U485  ( .a(\comparator/N1560 ), .out(\comparator/n485 ) );
  inv \comparator/U484  ( .a(\comparator/N1563 ), .out(\comparator/n484 ) );
  inv \comparator/U483  ( .a(\comparator/N1562 ), .out(\comparator/n483 ) );
  inv \comparator/U482  ( .a(\comparator/N1565 ), .out(\comparator/n482 ) );
  inv \comparator/U481  ( .a(\comparator/N1564 ), .out(\comparator/n481 ) );
  inv \comparator/U480  ( .a(\comparator/N1567 ), .out(\comparator/n480 ) );
  inv \comparator/U479  ( .a(\comparator/N1566 ), .out(\comparator/n479 ) );
  inv \comparator/U478  ( .a(\comparator/N1569 ), .out(\comparator/n478 ) );
  inv \comparator/U477  ( .a(\comparator/N1568 ), .out(\comparator/n477 ) );
  inv \comparator/U476  ( .a(\comparator/N1571 ), .out(\comparator/n476 ) );
  inv \comparator/U475  ( .a(\comparator/N1570 ), .out(\comparator/n475 ) );
  inv \comparator/U474  ( .a(\comparator/N1573 ), .out(\comparator/n474 ) );
  inv \comparator/U473  ( .a(\comparator/N1572 ), .out(\comparator/n473 ) );
  inv \comparator/U472  ( .a(\comparator/N1575 ), .out(\comparator/n472 ) );
  inv \comparator/U471  ( .a(\comparator/N1574 ), .out(\comparator/n471 ) );
  inv \comparator/U470  ( .a(\comparator/N1577 ), .out(\comparator/n470 ) );
  inv \comparator/U469  ( .a(\comparator/N1576 ), .out(\comparator/n469 ) );
  inv \comparator/U468  ( .a(\comparator/N1579 ), .out(\comparator/n468 ) );
  inv \comparator/U467  ( .a(\comparator/N1578 ), .out(\comparator/n467 ) );
  inv \comparator/U466  ( .a(\comparator/N1581 ), .out(\comparator/n466 ) );
  inv \comparator/U465  ( .a(\comparator/N1580 ), .out(\comparator/n465 ) );
  inv \comparator/U464  ( .a(\comparator/N1583 ), .out(\comparator/n464 ) );
  inv \comparator/U463  ( .a(\comparator/N1582 ), .out(\comparator/n463 ) );
  inv \comparator/U462  ( .a(\comparator/N1585 ), .out(\comparator/n462 ) );
  inv \comparator/U461  ( .a(\comparator/N1584 ), .out(\comparator/n461 ) );
  inv \comparator/U460  ( .a(\comparator/N1587 ), .out(\comparator/n460 ) );
  inv \comparator/U459  ( .a(\comparator/N1586 ), .out(\comparator/n459 ) );
  inv \comparator/U458  ( .a(\comparator/N1589 ), .out(\comparator/n458 ) );
  inv \comparator/U457  ( .a(\comparator/N1588 ), .out(\comparator/n457 ) );
  inv \comparator/U456  ( .a(\comparator/N1591 ), .out(\comparator/n456 ) );
  inv \comparator/U455  ( .a(\comparator/N1590 ), .out(\comparator/n455 ) );
  inv \comparator/U454  ( .a(\comparator/N1593 ), .out(\comparator/n454 ) );
  inv \comparator/U453  ( .a(\comparator/N1592 ), .out(\comparator/n453 ) );
  inv \comparator/U452  ( .a(\comparator/N1595 ), .out(\comparator/n452 ) );
  inv \comparator/U451  ( .a(\comparator/N1594 ), .out(\comparator/n451 ) );
  inv \comparator/U450  ( .a(\comparator/N1597 ), .out(\comparator/n450 ) );
  inv \comparator/U449  ( .a(\comparator/N1596 ), .out(\comparator/n449 ) );
  inv \comparator/U448  ( .a(\comparator/N1599 ), .out(\comparator/n448 ) );
  inv \comparator/U447  ( .a(\comparator/N1598 ), .out(\comparator/n447 ) );
  inv \comparator/U446  ( .a(\comparator/N1601 ), .out(\comparator/n446 ) );
  inv \comparator/U445  ( .a(\comparator/N1600 ), .out(\comparator/n445 ) );
  inv \comparator/U444  ( .a(\comparator/N1603 ), .out(\comparator/n444 ) );
  inv \comparator/U443  ( .a(\comparator/N1602 ), .out(\comparator/n443 ) );
  inv \comparator/U442  ( .a(\comparator/N1605 ), .out(\comparator/n442 ) );
  inv \comparator/U441  ( .a(\comparator/N1604 ), .out(\comparator/n441 ) );
  inv \comparator/U440  ( .a(\comparator/N1607 ), .out(\comparator/n440 ) );
  inv \comparator/U439  ( .a(\comparator/N1606 ), .out(\comparator/n439 ) );
  inv \comparator/U438  ( .a(\comparator/N1609 ), .out(\comparator/n438 ) );
  inv \comparator/U437  ( .a(\comparator/N1608 ), .out(\comparator/n437 ) );
  inv \comparator/U436  ( .a(\comparator/N1611 ), .out(\comparator/n436 ) );
  inv \comparator/U435  ( .a(\comparator/N1610 ), .out(\comparator/n435 ) );
  inv \comparator/U434  ( .a(\comparator/N1613 ), .out(\comparator/n434 ) );
  inv \comparator/U433  ( .a(\comparator/N1612 ), .out(\comparator/n433 ) );
  inv \comparator/U432  ( .a(\comparator/N1615 ), .out(\comparator/n432 ) );
  inv \comparator/U431  ( .a(\comparator/N1614 ), .out(\comparator/n431 ) );
  inv \comparator/U430  ( .a(\comparator/N1617 ), .out(\comparator/n430 ) );
  inv \comparator/U429  ( .a(\comparator/N1616 ), .out(\comparator/n429 ) );
  inv \comparator/U428  ( .a(\comparator/N1619 ), .out(\comparator/n428 ) );
  inv \comparator/U427  ( .a(\comparator/N1618 ), .out(\comparator/n427 ) );
  inv \comparator/U426  ( .a(\comparator/N1621 ), .out(\comparator/n426 ) );
  inv \comparator/U425  ( .a(\comparator/N1620 ), .out(\comparator/n425 ) );
  inv \comparator/U424  ( .a(\comparator/N1623 ), .out(\comparator/n424 ) );
  inv \comparator/U423  ( .a(\comparator/N1622 ), .out(\comparator/n423 ) );
  inv \comparator/U422  ( .a(\comparator/N1625 ), .out(\comparator/n422 ) );
  inv \comparator/U421  ( .a(\comparator/N1624 ), .out(\comparator/n421 ) );
  inv \comparator/U420  ( .a(\comparator/N1627 ), .out(\comparator/n420 ) );
  inv \comparator/U419  ( .a(\comparator/N1626 ), .out(\comparator/n419 ) );
  inv \comparator/U418  ( .a(\comparator/N1629 ), .out(\comparator/n418 ) );
  inv \comparator/U417  ( .a(\comparator/N1628 ), .out(\comparator/n417 ) );
  inv \comparator/U416  ( .a(\comparator/N1631 ), .out(\comparator/n416 ) );
  inv \comparator/U415  ( .a(\comparator/N1630 ), .out(\comparator/n415 ) );
  inv \comparator/U414  ( .a(\comparator/N1633 ), .out(\comparator/n414 ) );
  inv \comparator/U413  ( .a(\comparator/N1632 ), .out(\comparator/n413 ) );
  inv \comparator/U412  ( .a(\comparator/N1635 ), .out(\comparator/n412 ) );
  inv \comparator/U411  ( .a(\comparator/N1634 ), .out(\comparator/n411 ) );
  inv \comparator/U410  ( .a(\comparator/N1637 ), .out(\comparator/n410 ) );
  inv \comparator/U409  ( .a(\comparator/N1636 ), .out(\comparator/n409 ) );
  inv \comparator/U408  ( .a(\comparator/N1639 ), .out(\comparator/n408 ) );
  inv \comparator/U407  ( .a(\comparator/N1638 ), .out(\comparator/n407 ) );
  inv \comparator/U406  ( .a(\comparator/N1641 ), .out(\comparator/n406 ) );
  inv \comparator/U405  ( .a(\comparator/N1640 ), .out(\comparator/n405 ) );
  inv \comparator/U404  ( .a(\comparator/N1643 ), .out(\comparator/n404 ) );
  inv \comparator/U403  ( .a(\comparator/N1642 ), .out(\comparator/n403 ) );
  inv \comparator/U402  ( .a(\comparator/N1645 ), .out(\comparator/n402 ) );
  inv \comparator/U401  ( .a(\comparator/N1644 ), .out(\comparator/n401 ) );
  inv \comparator/U400  ( .a(\comparator/N1647 ), .out(\comparator/n400 ) );
  inv \comparator/U399  ( .a(\comparator/N1646 ), .out(\comparator/n399 ) );
  inv \comparator/U398  ( .a(\comparator/N1649 ), .out(\comparator/n398 ) );
  inv \comparator/U397  ( .a(\comparator/N1648 ), .out(\comparator/n397 ) );
  inv \comparator/U396  ( .a(\comparator/N1651 ), .out(\comparator/n396 ) );
  inv \comparator/U395  ( .a(\comparator/N1650 ), .out(\comparator/n395 ) );
  inv \comparator/U394  ( .a(\comparator/N1653 ), .out(\comparator/n394 ) );
  inv \comparator/U393  ( .a(\comparator/N1652 ), .out(\comparator/n393 ) );
  inv \comparator/U392  ( .a(\comparator/N1655 ), .out(\comparator/n392 ) );
  inv \comparator/U391  ( .a(\comparator/N1654 ), .out(\comparator/n391 ) );
  inv \comparator/U390  ( .a(\comparator/N1657 ), .out(\comparator/n390 ) );
  inv \comparator/U389  ( .a(\comparator/N1656 ), .out(\comparator/n389 ) );
  inv \comparator/U388  ( .a(\comparator/N1659 ), .out(\comparator/n388 ) );
  inv \comparator/U387  ( .a(\comparator/N1658 ), .out(\comparator/n387 ) );
  inv \comparator/U386  ( .a(\comparator/N1661 ), .out(\comparator/n386 ) );
  inv \comparator/U385  ( .a(\comparator/N1660 ), .out(\comparator/n385 ) );
  inv \comparator/U384  ( .a(\comparator/N1663 ), .out(\comparator/n384 ) );
  inv \comparator/U383  ( .a(\comparator/N1662 ), .out(\comparator/n383 ) );
  inv \comparator/U382  ( .a(\comparator/N1665 ), .out(\comparator/n382 ) );
  inv \comparator/U381  ( .a(\comparator/N1664 ), .out(\comparator/n381 ) );
  inv \comparator/U380  ( .a(\comparator/N1667 ), .out(\comparator/n380 ) );
  inv \comparator/U379  ( .a(\comparator/N1666 ), .out(\comparator/n379 ) );
  inv \comparator/U378  ( .a(\comparator/N1669 ), .out(\comparator/n378 ) );
  inv \comparator/U377  ( .a(\comparator/N1668 ), .out(\comparator/n377 ) );
  inv \comparator/U376  ( .a(\comparator/N1671 ), .out(\comparator/n376 ) );
  inv \comparator/U375  ( .a(\comparator/N1670 ), .out(\comparator/n375 ) );
  inv \comparator/U374  ( .a(\comparator/N1673 ), .out(\comparator/n374 ) );
  inv \comparator/U373  ( .a(\comparator/N1672 ), .out(\comparator/n373 ) );
  inv \comparator/U372  ( .a(\comparator/N1675 ), .out(\comparator/n372 ) );
  inv \comparator/U371  ( .a(\comparator/N1674 ), .out(\comparator/n371 ) );
  inv \comparator/U370  ( .a(\comparator/N1677 ), .out(\comparator/n370 ) );
  inv \comparator/U369  ( .a(\comparator/N1676 ), .out(\comparator/n369 ) );
  inv \comparator/U368  ( .a(\comparator/N1679 ), .out(\comparator/n368 ) );
  inv \comparator/U367  ( .a(\comparator/N1678 ), .out(\comparator/n367 ) );
  inv \comparator/U366  ( .a(\comparator/N1681 ), .out(\comparator/n366 ) );
  inv \comparator/U365  ( .a(\comparator/N1680 ), .out(\comparator/n365 ) );
  inv \comparator/U364  ( .a(\comparator/N1683 ), .out(\comparator/n364 ) );
  inv \comparator/U363  ( .a(\comparator/N1682 ), .out(\comparator/n363 ) );
  inv \comparator/U362  ( .a(\comparator/N1685 ), .out(\comparator/n362 ) );
  inv \comparator/U361  ( .a(\comparator/N1684 ), .out(\comparator/n361 ) );
  inv \comparator/U360  ( .a(\comparator/N1687 ), .out(\comparator/n360 ) );
  inv \comparator/U359  ( .a(\comparator/N1686 ), .out(\comparator/n359 ) );
  inv \comparator/U358  ( .a(\comparator/N1689 ), .out(\comparator/n358 ) );
  inv \comparator/U357  ( .a(\comparator/N1688 ), .out(\comparator/n357 ) );
  inv \comparator/U356  ( .a(\comparator/N1691 ), .out(\comparator/n356 ) );
  inv \comparator/U355  ( .a(\comparator/N1690 ), .out(\comparator/n355 ) );
  inv \comparator/U354  ( .a(\comparator/N1693 ), .out(\comparator/n354 ) );
  inv \comparator/U353  ( .a(\comparator/N1692 ), .out(\comparator/n353 ) );
  inv \comparator/U352  ( .a(\comparator/N1695 ), .out(\comparator/n352 ) );
  inv \comparator/U351  ( .a(\comparator/N1694 ), .out(\comparator/n351 ) );
  inv \comparator/U350  ( .a(\comparator/N1697 ), .out(\comparator/n350 ) );
  inv \comparator/U349  ( .a(\comparator/N1696 ), .out(\comparator/n349 ) );
  inv \comparator/U348  ( .a(\comparator/N1699 ), .out(\comparator/n348 ) );
  inv \comparator/U347  ( .a(\comparator/N1698 ), .out(\comparator/n347 ) );
  inv \comparator/U346  ( .a(\comparator/N1701 ), .out(\comparator/n346 ) );
  inv \comparator/U345  ( .a(\comparator/N1700 ), .out(\comparator/n345 ) );
  inv \comparator/U344  ( .a(\comparator/N1703 ), .out(\comparator/n344 ) );
  inv \comparator/U343  ( .a(\comparator/N1702 ), .out(\comparator/n343 ) );
  inv \comparator/U342  ( .a(\comparator/N1705 ), .out(\comparator/n342 ) );
  inv \comparator/U341  ( .a(\comparator/N1704 ), .out(\comparator/n341 ) );
  inv \comparator/U340  ( .a(\comparator/N1707 ), .out(\comparator/n340 ) );
  inv \comparator/U339  ( .a(\comparator/N1706 ), .out(\comparator/n339 ) );
  inv \comparator/U338  ( .a(\comparator/N1709 ), .out(\comparator/n338 ) );
  inv \comparator/U337  ( .a(\comparator/N1708 ), .out(\comparator/n337 ) );
  inv \comparator/U336  ( .a(\comparator/N1711 ), .out(\comparator/n336 ) );
  inv \comparator/U335  ( .a(\comparator/N1710 ), .out(\comparator/n335 ) );
  inv \comparator/U334  ( .a(\comparator/N1713 ), .out(\comparator/n334 ) );
  inv \comparator/U333  ( .a(\comparator/N1712 ), .out(\comparator/n333 ) );
  inv \comparator/U332  ( .a(\comparator/N1715 ), .out(\comparator/n332 ) );
  inv \comparator/U331  ( .a(\comparator/N1714 ), .out(\comparator/n331 ) );
  inv \comparator/U330  ( .a(\comparator/N1717 ), .out(\comparator/n330 ) );
  inv \comparator/U329  ( .a(\comparator/N1716 ), .out(\comparator/n329 ) );
  inv \comparator/U328  ( .a(\comparator/N1719 ), .out(\comparator/n328 ) );
  inv \comparator/U327  ( .a(\comparator/N1718 ), .out(\comparator/n327 ) );
  inv \comparator/U326  ( .a(\comparator/N1721 ), .out(\comparator/n326 ) );
  inv \comparator/U325  ( .a(\comparator/N1720 ), .out(\comparator/n325 ) );
  inv \comparator/U324  ( .a(\comparator/N1723 ), .out(\comparator/n324 ) );
  inv \comparator/U323  ( .a(\comparator/N1722 ), .out(\comparator/n323 ) );
  inv \comparator/U322  ( .a(\comparator/N1725 ), .out(\comparator/n322 ) );
  inv \comparator/U321  ( .a(\comparator/N1724 ), .out(\comparator/n321 ) );
  inv \comparator/U320  ( .a(\comparator/N1727 ), .out(\comparator/n320 ) );
  inv \comparator/U319  ( .a(\comparator/N1726 ), .out(\comparator/n319 ) );
  inv \comparator/U318  ( .a(\comparator/N1729 ), .out(\comparator/n318 ) );
  inv \comparator/U317  ( .a(\comparator/N1728 ), .out(\comparator/n317 ) );
  inv \comparator/U316  ( .a(\comparator/N1731 ), .out(\comparator/n316 ) );
  inv \comparator/U315  ( .a(\comparator/N1730 ), .out(\comparator/n315 ) );
  inv \comparator/U314  ( .a(\comparator/N1733 ), .out(\comparator/n314 ) );
  inv \comparator/U313  ( .a(\comparator/N1732 ), .out(\comparator/n313 ) );
  inv \comparator/U312  ( .a(\comparator/N1735 ), .out(\comparator/n312 ) );
  inv \comparator/U311  ( .a(\comparator/N1734 ), .out(\comparator/n311 ) );
  inv \comparator/U310  ( .a(\comparator/N1737 ), .out(\comparator/n310 ) );
  inv \comparator/U309  ( .a(\comparator/N1736 ), .out(\comparator/n309 ) );
  inv \comparator/U308  ( .a(\comparator/N1739 ), .out(\comparator/n308 ) );
  inv \comparator/U307  ( .a(\comparator/N1738 ), .out(\comparator/n307 ) );
  inv \comparator/U306  ( .a(\comparator/N1741 ), .out(\comparator/n306 ) );
  inv \comparator/U305  ( .a(\comparator/N1740 ), .out(\comparator/n305 ) );
  inv \comparator/U304  ( .a(\comparator/N1743 ), .out(\comparator/n304 ) );
  inv \comparator/U303  ( .a(\comparator/N1742 ), .out(\comparator/n303 ) );
  inv \comparator/U302  ( .a(\comparator/N1745 ), .out(\comparator/n302 ) );
  inv \comparator/U301  ( .a(\comparator/N1744 ), .out(\comparator/n301 ) );
  inv \comparator/U300  ( .a(\comparator/N1747 ), .out(\comparator/n300 ) );
  inv \comparator/U299  ( .a(\comparator/N1746 ), .out(\comparator/n299 ) );
  inv \comparator/U298  ( .a(\comparator/N1749 ), .out(\comparator/n298 ) );
  inv \comparator/U297  ( .a(\comparator/N1748 ), .out(\comparator/n297 ) );
  inv \comparator/U296  ( .a(\comparator/N1751 ), .out(\comparator/n296 ) );
  inv \comparator/U295  ( .a(\comparator/N1750 ), .out(\comparator/n295 ) );
  inv \comparator/U294  ( .a(\comparator/N1753 ), .out(\comparator/n294 ) );
  inv \comparator/U293  ( .a(\comparator/N1752 ), .out(\comparator/n293 ) );
  inv \comparator/U292  ( .a(\comparator/N1755 ), .out(\comparator/n292 ) );
  inv \comparator/U291  ( .a(\comparator/N1754 ), .out(\comparator/n291 ) );
  inv \comparator/U290  ( .a(\comparator/N1757 ), .out(\comparator/n290 ) );
  inv \comparator/U289  ( .a(\comparator/N1756 ), .out(\comparator/n289 ) );
  inv \comparator/U288  ( .a(\comparator/N1759 ), .out(\comparator/n288 ) );
  inv \comparator/U287  ( .a(\comparator/N1758 ), .out(\comparator/n287 ) );
  inv \comparator/U286  ( .a(\comparator/N1761 ), .out(\comparator/n286 ) );
  inv \comparator/U285  ( .a(\comparator/N1760 ), .out(\comparator/n285 ) );
  inv \comparator/U284  ( .a(\comparator/N1763 ), .out(\comparator/n284 ) );
  inv \comparator/U283  ( .a(\comparator/N1762 ), .out(\comparator/n283 ) );
  inv \comparator/U282  ( .a(\comparator/N1765 ), .out(\comparator/n282 ) );
  inv \comparator/U281  ( .a(\comparator/N1764 ), .out(\comparator/n281 ) );
  inv \comparator/U280  ( .a(\comparator/N1767 ), .out(\comparator/n280 ) );
  inv \comparator/U279  ( .a(\comparator/N1766 ), .out(\comparator/n279 ) );
  inv \comparator/U278  ( .a(\comparator/N1769 ), .out(\comparator/n278 ) );
  inv \comparator/U277  ( .a(\comparator/N1768 ), .out(\comparator/n277 ) );
  inv \comparator/U276  ( .a(\comparator/N1771 ), .out(\comparator/n276 ) );
  inv \comparator/U275  ( .a(\comparator/N1770 ), .out(\comparator/n275 ) );
  inv \comparator/U274  ( .a(\comparator/N1773 ), .out(\comparator/n274 ) );
  inv \comparator/U273  ( .a(\comparator/N1772 ), .out(\comparator/n273 ) );
  inv \comparator/U272  ( .a(\comparator/N1775 ), .out(\comparator/n272 ) );
  inv \comparator/U271  ( .a(\comparator/N1774 ), .out(\comparator/n271 ) );
  inv \comparator/U270  ( .a(\comparator/N1777 ), .out(\comparator/n270 ) );
  inv \comparator/U269  ( .a(\comparator/N1776 ), .out(\comparator/n269 ) );
  inv \comparator/U268  ( .a(\comparator/N1779 ), .out(\comparator/n268 ) );
  inv \comparator/U267  ( .a(\comparator/N1778 ), .out(\comparator/n267 ) );
  inv \comparator/U266  ( .a(\comparator/N1781 ), .out(\comparator/n266 ) );
  inv \comparator/U265  ( .a(\comparator/N1780 ), .out(\comparator/n265 ) );
  inv \comparator/U264  ( .a(\comparator/N1783 ), .out(\comparator/n264 ) );
  inv \comparator/U263  ( .a(\comparator/N1782 ), .out(\comparator/n263 ) );
  inv \comparator/U262  ( .a(\comparator/N1785 ), .out(\comparator/n262 ) );
  inv \comparator/U261  ( .a(\comparator/N1784 ), .out(\comparator/n261 ) );
  inv \comparator/U260  ( .a(\comparator/N1787 ), .out(\comparator/n260 ) );
  inv \comparator/U259  ( .a(\comparator/N1786 ), .out(\comparator/n259 ) );
  inv \comparator/U258  ( .a(\comparator/N1789 ), .out(\comparator/n258 ) );
  inv \comparator/U257  ( .a(\comparator/N1788 ), .out(\comparator/n257 ) );
  inv \comparator/U256  ( .a(\comparator/N1791 ), .out(\comparator/n256 ) );
  inv \comparator/U255  ( .a(\comparator/N1790 ), .out(\comparator/n255 ) );
  inv \comparator/U254  ( .a(\comparator/N1793 ), .out(\comparator/n254 ) );
  inv \comparator/U253  ( .a(\comparator/N1792 ), .out(\comparator/n253 ) );
  inv \comparator/U252  ( .a(\comparator/N1795 ), .out(\comparator/n252 ) );
  inv \comparator/U251  ( .a(\comparator/N1794 ), .out(\comparator/n251 ) );
  inv \comparator/U250  ( .a(\comparator/N1797 ), .out(\comparator/n250 ) );
  inv \comparator/U249  ( .a(\comparator/N1796 ), .out(\comparator/n249 ) );
  inv \comparator/U248  ( .a(\comparator/N1799 ), .out(\comparator/n248 ) );
  inv \comparator/U247  ( .a(\comparator/N1798 ), .out(\comparator/n247 ) );
  inv \comparator/U246  ( .a(\comparator/N1801 ), .out(\comparator/n246 ) );
  inv \comparator/U245  ( .a(\comparator/N1800 ), .out(\comparator/n245 ) );
  inv \comparator/U244  ( .a(\comparator/N1803 ), .out(\comparator/n244 ) );
  inv \comparator/U243  ( .a(\comparator/N1802 ), .out(\comparator/n243 ) );
  inv \comparator/U242  ( .a(\comparator/N1805 ), .out(\comparator/n242 ) );
  inv \comparator/U241  ( .a(\comparator/N1804 ), .out(\comparator/n241 ) );
  inv \comparator/U240  ( .a(\comparator/N1807 ), .out(\comparator/n240 ) );
  inv \comparator/U239  ( .a(\comparator/N1806 ), .out(\comparator/n239 ) );
  inv \comparator/U238  ( .a(\comparator/N1809 ), .out(\comparator/n238 ) );
  inv \comparator/U237  ( .a(\comparator/N1808 ), .out(\comparator/n237 ) );
  inv \comparator/U236  ( .a(\comparator/N1811 ), .out(\comparator/n236 ) );
  inv \comparator/U235  ( .a(\comparator/N1810 ), .out(\comparator/n235 ) );
  inv \comparator/U234  ( .a(\comparator/N1813 ), .out(\comparator/n234 ) );
  inv \comparator/U233  ( .a(\comparator/N1812 ), .out(\comparator/n233 ) );
  inv \comparator/U232  ( .a(\comparator/N1815 ), .out(\comparator/n232 ) );
  inv \comparator/U231  ( .a(\comparator/N1814 ), .out(\comparator/n231 ) );
  inv \comparator/U230  ( .a(\comparator/N1817 ), .out(\comparator/n230 ) );
  inv \comparator/U229  ( .a(\comparator/N1816 ), .out(\comparator/n229 ) );
  inv \comparator/U228  ( .a(\comparator/N1819 ), .out(\comparator/n228 ) );
  inv \comparator/U227  ( .a(\comparator/N1818 ), .out(\comparator/n227 ) );
  inv \comparator/U226  ( .a(\comparator/N1821 ), .out(\comparator/n226 ) );
  inv \comparator/U225  ( .a(\comparator/N1820 ), .out(\comparator/n225 ) );
  inv \comparator/U224  ( .a(\comparator/N1823 ), .out(\comparator/n224 ) );
  inv \comparator/U223  ( .a(\comparator/N1822 ), .out(\comparator/n223 ) );
  inv \comparator/U222  ( .a(\comparator/N1825 ), .out(\comparator/n222 ) );
  inv \comparator/U221  ( .a(\comparator/N1824 ), .out(\comparator/n221 ) );
  inv \comparator/U220  ( .a(\comparator/N1827 ), .out(\comparator/n220 ) );
  inv \comparator/U219  ( .a(\comparator/N1826 ), .out(\comparator/n219 ) );
  inv \comparator/U218  ( .a(\comparator/N1829 ), .out(\comparator/n218 ) );
  inv \comparator/U217  ( .a(\comparator/N1828 ), .out(\comparator/n217 ) );
  inv \comparator/U216  ( .a(\comparator/N1831 ), .out(\comparator/n216 ) );
  inv \comparator/U215  ( .a(\comparator/N1830 ), .out(\comparator/n215 ) );
  inv \comparator/U214  ( .a(\comparator/N1833 ), .out(\comparator/n214 ) );
  inv \comparator/U213  ( .a(\comparator/N1832 ), .out(\comparator/n213 ) );
  inv \comparator/U212  ( .a(\comparator/N1835 ), .out(\comparator/n212 ) );
  inv \comparator/U211  ( .a(\comparator/N1834 ), .out(\comparator/n211 ) );
  inv \comparator/U210  ( .a(\comparator/N1837 ), .out(\comparator/n210 ) );
  inv \comparator/U209  ( .a(\comparator/N1836 ), .out(\comparator/n209 ) );
  inv \comparator/U208  ( .a(\comparator/N1839 ), .out(\comparator/n208 ) );
  inv \comparator/U207  ( .a(\comparator/N1838 ), .out(\comparator/n207 ) );
  inv \comparator/U206  ( .a(\comparator/N1841 ), .out(\comparator/n206 ) );
  inv \comparator/U205  ( .a(\comparator/N1840 ), .out(\comparator/n205 ) );
  inv \comparator/U204  ( .a(\comparator/N1843 ), .out(\comparator/n204 ) );
  inv \comparator/U203  ( .a(\comparator/N1842 ), .out(\comparator/n203 ) );
  inv \comparator/U202  ( .a(\comparator/N1845 ), .out(\comparator/n202 ) );
  inv \comparator/U201  ( .a(\comparator/N1844 ), .out(\comparator/n201 ) );
  inv \comparator/U200  ( .a(\comparator/N1847 ), .out(\comparator/n200 ) );
  inv \comparator/U199  ( .a(\comparator/N1846 ), .out(\comparator/n199 ) );
  inv \comparator/U198  ( .a(\comparator/N1849 ), .out(\comparator/n198 ) );
  inv \comparator/U197  ( .a(\comparator/N1848 ), .out(\comparator/n197 ) );
  inv \comparator/U196  ( .a(\comparator/N1851 ), .out(\comparator/n196 ) );
  inv \comparator/U195  ( .a(\comparator/N1850 ), .out(\comparator/n195 ) );
  inv \comparator/U194  ( .a(\comparator/N1853 ), .out(\comparator/n194 ) );
  inv \comparator/U193  ( .a(\comparator/N1852 ), .out(\comparator/n193 ) );
  inv \comparator/U192  ( .a(\comparator/N1855 ), .out(\comparator/n192 ) );
  inv \comparator/U191  ( .a(\comparator/N1854 ), .out(\comparator/n191 ) );
  inv \comparator/U190  ( .a(\comparator/N1857 ), .out(\comparator/n190 ) );
  inv \comparator/U189  ( .a(\comparator/N1856 ), .out(\comparator/n189 ) );
  inv \comparator/U188  ( .a(\comparator/N1859 ), .out(\comparator/n188 ) );
  inv \comparator/U187  ( .a(\comparator/N1858 ), .out(\comparator/n187 ) );
  inv \comparator/U186  ( .a(\comparator/N1861 ), .out(\comparator/n186 ) );
  inv \comparator/U185  ( .a(\comparator/N1860 ), .out(\comparator/n185 ) );
  inv \comparator/U184  ( .a(\comparator/N1863 ), .out(\comparator/n184 ) );
  inv \comparator/U183  ( .a(\comparator/N1862 ), .out(\comparator/n183 ) );
  inv \comparator/U182  ( .a(\comparator/N1865 ), .out(\comparator/n182 ) );
  inv \comparator/U181  ( .a(\comparator/N1864 ), .out(\comparator/n181 ) );
  inv \comparator/U180  ( .a(\comparator/N1867 ), .out(\comparator/n180 ) );
  inv \comparator/U179  ( .a(\comparator/N1866 ), .out(\comparator/n179 ) );
  inv \comparator/U178  ( .a(\comparator/N1869 ), .out(\comparator/n178 ) );
  inv \comparator/U177  ( .a(\comparator/N1868 ), .out(\comparator/n177 ) );
  inv \comparator/U176  ( .a(\comparator/N1871 ), .out(\comparator/n176 ) );
  inv \comparator/U175  ( .a(\comparator/N1870 ), .out(\comparator/n175 ) );
  inv \comparator/U174  ( .a(\comparator/N1873 ), .out(\comparator/n174 ) );
  inv \comparator/U173  ( .a(\comparator/N1872 ), .out(\comparator/n173 ) );
  inv \comparator/U172  ( .a(\comparator/N1875 ), .out(\comparator/n172 ) );
  inv \comparator/U171  ( .a(\comparator/N1874 ), .out(\comparator/n171 ) );
  inv \comparator/U170  ( .a(\comparator/N1877 ), .out(\comparator/n170 ) );
  inv \comparator/U169  ( .a(\comparator/N1876 ), .out(\comparator/n169 ) );
  inv \comparator/U168  ( .a(\comparator/N1879 ), .out(\comparator/n168 ) );
  inv \comparator/U167  ( .a(\comparator/N1878 ), .out(\comparator/n167 ) );
  inv \comparator/U166  ( .a(\comparator/N1881 ), .out(\comparator/n166 ) );
  inv \comparator/U165  ( .a(\comparator/N1880 ), .out(\comparator/n165 ) );
  inv \comparator/U164  ( .a(\comparator/N1883 ), .out(\comparator/n164 ) );
  inv \comparator/U163  ( .a(\comparator/N1882 ), .out(\comparator/n163 ) );
  inv \comparator/U162  ( .a(\comparator/N1885 ), .out(\comparator/n162 ) );
  inv \comparator/U161  ( .a(\comparator/N1884 ), .out(\comparator/n161 ) );
  inv \comparator/U160  ( .a(\comparator/N1887 ), .out(\comparator/n160 ) );
  inv \comparator/U159  ( .a(\comparator/N1886 ), .out(\comparator/n159 ) );
  inv \comparator/U158  ( .a(\comparator/N1889 ), .out(\comparator/n158 ) );
  inv \comparator/U157  ( .a(\comparator/N1888 ), .out(\comparator/n157 ) );
  inv \comparator/U156  ( .a(\comparator/N1891 ), .out(\comparator/n156 ) );
  inv \comparator/U155  ( .a(\comparator/N1890 ), .out(\comparator/n155 ) );
  inv \comparator/U154  ( .a(\comparator/N1893 ), .out(\comparator/n154 ) );
  inv \comparator/U153  ( .a(\comparator/N1892 ), .out(\comparator/n153 ) );
  inv \comparator/U152  ( .a(\comparator/N1895 ), .out(\comparator/n152 ) );
  inv \comparator/U151  ( .a(\comparator/N1894 ), .out(\comparator/n151 ) );
  inv \comparator/U150  ( .a(\comparator/N1897 ), .out(\comparator/n150 ) );
  inv \comparator/U149  ( .a(\comparator/N1896 ), .out(\comparator/n149 ) );
  inv \comparator/U148  ( .a(\comparator/N1899 ), .out(\comparator/n148 ) );
  inv \comparator/U147  ( .a(\comparator/N1898 ), .out(\comparator/n147 ) );
  inv \comparator/U146  ( .a(\comparator/N1901 ), .out(\comparator/n146 ) );
  inv \comparator/U145  ( .a(\comparator/N1900 ), .out(\comparator/n145 ) );
  inv \comparator/U144  ( .a(\comparator/N1903 ), .out(\comparator/n144 ) );
  inv \comparator/U143  ( .a(\comparator/N1902 ), .out(\comparator/n143 ) );
  inv \comparator/U142  ( .a(\comparator/N1905 ), .out(\comparator/n142 ) );
  inv \comparator/U141  ( .a(\comparator/N1904 ), .out(\comparator/n141 ) );
  inv \comparator/U140  ( .a(\comparator/N1907 ), .out(\comparator/n140 ) );
  inv \comparator/U139  ( .a(\comparator/N1906 ), .out(\comparator/n139 ) );
  inv \comparator/U138  ( .a(\comparator/N1909 ), .out(\comparator/n138 ) );
  inv \comparator/U137  ( .a(\comparator/N1908 ), .out(\comparator/n137 ) );
  inv \comparator/U136  ( .a(\comparator/N1911 ), .out(\comparator/n136 ) );
  inv \comparator/U135  ( .a(\comparator/N1910 ), .out(\comparator/n135 ) );
  inv \comparator/U134  ( .a(\comparator/N1913 ), .out(\comparator/n134 ) );
  inv \comparator/U133  ( .a(\comparator/N1912 ), .out(\comparator/n133 ) );
  inv \comparator/U132  ( .a(\comparator/N1915 ), .out(\comparator/n132 ) );
  inv \comparator/U131  ( .a(\comparator/N1914 ), .out(\comparator/n131 ) );
  inv \comparator/U130  ( .a(\comparator/N1917 ), .out(\comparator/n130 ) );
  inv \comparator/U129  ( .a(\comparator/N1916 ), .out(\comparator/n129 ) );
  inv \comparator/U128  ( .a(\comparator/N1919 ), .out(\comparator/n128 ) );
  inv \comparator/U127  ( .a(\comparator/N1918 ), .out(\comparator/n127 ) );
  inv \comparator/U126  ( .a(\comparator/N1921 ), .out(\comparator/n126 ) );
  inv \comparator/U125  ( .a(\comparator/N1920 ), .out(\comparator/n125 ) );
  inv \comparator/U124  ( .a(\comparator/N1923 ), .out(\comparator/n124 ) );
  inv \comparator/U123  ( .a(\comparator/N1922 ), .out(\comparator/n123 ) );
  inv \comparator/U122  ( .a(\comparator/N1925 ), .out(\comparator/n122 ) );
  inv \comparator/U121  ( .a(\comparator/N1924 ), .out(\comparator/n121 ) );
  inv \comparator/U120  ( .a(\comparator/N1927 ), .out(\comparator/n120 ) );
  inv \comparator/U119  ( .a(\comparator/N1926 ), .out(\comparator/n119 ) );
  inv \comparator/U118  ( .a(\comparator/N1929 ), .out(\comparator/n118 ) );
  inv \comparator/U117  ( .a(\comparator/N1928 ), .out(\comparator/n117 ) );
  inv \comparator/U116  ( .a(\comparator/N1931 ), .out(\comparator/n116 ) );
  inv \comparator/U115  ( .a(\comparator/N1930 ), .out(\comparator/n115 ) );
  inv \comparator/U114  ( .a(\comparator/N1933 ), .out(\comparator/n114 ) );
  inv \comparator/U113  ( .a(\comparator/N1932 ), .out(\comparator/n113 ) );
  inv \comparator/U112  ( .a(\comparator/N1935 ), .out(\comparator/n112 ) );
  inv \comparator/U111  ( .a(\comparator/N1934 ), .out(\comparator/n111 ) );
  inv \comparator/U110  ( .a(\comparator/N1937 ), .out(\comparator/n110 ) );
  inv \comparator/U109  ( .a(\comparator/N1936 ), .out(\comparator/n109 ) );
  inv \comparator/U108  ( .a(\comparator/N1939 ), .out(\comparator/n108 ) );
  inv \comparator/U107  ( .a(\comparator/N1938 ), .out(\comparator/n107 ) );
  inv \comparator/U106  ( .a(\comparator/N1941 ), .out(\comparator/n106 ) );
  inv \comparator/U105  ( .a(\comparator/N1940 ), .out(\comparator/n105 ) );
  inv \comparator/U104  ( .a(\comparator/N1943 ), .out(\comparator/n104 ) );
  inv \comparator/U103  ( .a(\comparator/N1942 ), .out(\comparator/n103 ) );
  inv \comparator/U102  ( .a(\comparator/N1945 ), .out(\comparator/n102 ) );
  inv \comparator/U101  ( .a(\comparator/N1944 ), .out(\comparator/n101 ) );
  inv \comparator/U100  ( .a(\comparator/N1947 ), .out(\comparator/n100 ) );
  inv \comparator/U99  ( .a(\comparator/N1946 ), .out(\comparator/n99 ) );
  inv \comparator/U98  ( .a(\comparator/N1949 ), .out(\comparator/n98 ) );
  inv \comparator/U97  ( .a(\comparator/N1948 ), .out(\comparator/n97 ) );
  inv \comparator/U96  ( .a(\comparator/N1951 ), .out(\comparator/n96 ) );
  inv \comparator/U95  ( .a(\comparator/N1950 ), .out(\comparator/n95 ) );
  inv \comparator/U94  ( .a(\comparator/N1953 ), .out(\comparator/n94 ) );
  inv \comparator/U93  ( .a(\comparator/N1952 ), .out(\comparator/n93 ) );
  inv \comparator/U92  ( .a(\comparator/N1955 ), .out(\comparator/n92 ) );
  inv \comparator/U91  ( .a(\comparator/N1954 ), .out(\comparator/n91 ) );
  inv \comparator/U90  ( .a(\comparator/N1957 ), .out(\comparator/n90 ) );
  inv \comparator/U89  ( .a(\comparator/N1956 ), .out(\comparator/n89 ) );
  inv \comparator/U88  ( .a(\comparator/N1959 ), .out(\comparator/n88 ) );
  inv \comparator/U87  ( .a(\comparator/N1958 ), .out(\comparator/n87 ) );
  inv \comparator/U86  ( .a(\comparator/N1961 ), .out(\comparator/n86 ) );
  inv \comparator/U85  ( .a(\comparator/N1960 ), .out(\comparator/n85 ) );
  inv \comparator/U84  ( .a(\comparator/N1963 ), .out(\comparator/n84 ) );
  inv \comparator/U83  ( .a(\comparator/N1962 ), .out(\comparator/n83 ) );
  inv \comparator/U82  ( .a(\comparator/N1965 ), .out(\comparator/n82 ) );
  inv \comparator/U81  ( .a(\comparator/N1964 ), .out(\comparator/n81 ) );
  inv \comparator/U80  ( .a(\comparator/N1967 ), .out(\comparator/n80 ) );
  inv \comparator/U79  ( .a(\comparator/N1966 ), .out(\comparator/n79 ) );
  inv \comparator/U78  ( .a(\comparator/N1969 ), .out(\comparator/n78 ) );
  inv \comparator/U77  ( .a(\comparator/N1968 ), .out(\comparator/n77 ) );
  inv \comparator/U76  ( .a(\comparator/N1971 ), .out(\comparator/n76 ) );
  inv \comparator/U75  ( .a(\comparator/N1970 ), .out(\comparator/n75 ) );
  inv \comparator/U74  ( .a(\comparator/N1973 ), .out(\comparator/n74 ) );
  inv \comparator/U73  ( .a(\comparator/N1972 ), .out(\comparator/n73 ) );
  inv \comparator/U72  ( .a(\comparator/N1975 ), .out(\comparator/n72 ) );
  inv \comparator/U71  ( .a(\comparator/N1974 ), .out(\comparator/n71 ) );
  inv \comparator/U70  ( .a(\comparator/N1977 ), .out(\comparator/n70 ) );
  inv \comparator/U69  ( .a(\comparator/N1976 ), .out(\comparator/n69 ) );
  inv \comparator/U68  ( .a(\comparator/N1979 ), .out(\comparator/n68 ) );
  inv \comparator/U67  ( .a(\comparator/N1978 ), .out(\comparator/n67 ) );
  inv \comparator/U66  ( .a(\comparator/N1981 ), .out(\comparator/n66 ) );
  inv \comparator/U65  ( .a(\comparator/N1980 ), .out(\comparator/n65 ) );
  inv \comparator/U64  ( .a(\comparator/N1983 ), .out(\comparator/n64 ) );
  inv \comparator/U63  ( .a(\comparator/N1982 ), .out(\comparator/n63 ) );
  inv \comparator/U62  ( .a(\comparator/N1985 ), .out(\comparator/n62 ) );
  inv \comparator/U61  ( .a(\comparator/N1984 ), .out(\comparator/n61 ) );
  inv \comparator/U60  ( .a(\comparator/N1987 ), .out(\comparator/n60 ) );
  inv \comparator/U59  ( .a(\comparator/N1986 ), .out(\comparator/n59 ) );
  inv \comparator/U58  ( .a(\comparator/N1989 ), .out(\comparator/n58 ) );
  inv \comparator/U57  ( .a(\comparator/N1988 ), .out(\comparator/n57 ) );
  inv \comparator/U56  ( .a(\comparator/N1991 ), .out(\comparator/n56 ) );
  inv \comparator/U55  ( .a(\comparator/N1990 ), .out(\comparator/n55 ) );
  inv \comparator/U54  ( .a(\comparator/N1993 ), .out(\comparator/n54 ) );
  inv \comparator/U53  ( .a(\comparator/N1992 ), .out(\comparator/n53 ) );
  inv \comparator/U52  ( .a(\comparator/N1995 ), .out(\comparator/n52 ) );
  inv \comparator/U51  ( .a(\comparator/N1994 ), .out(\comparator/n51 ) );
  inv \comparator/U50  ( .a(\comparator/N1997 ), .out(\comparator/n50 ) );
  inv \comparator/U49  ( .a(\comparator/N1996 ), .out(\comparator/n49 ) );
  inv \comparator/U48  ( .a(\comparator/N1999 ), .out(\comparator/n48 ) );
  inv \comparator/U47  ( .a(\comparator/N1998 ), .out(\comparator/n47 ) );
  inv \comparator/U46  ( .a(\comparator/N2001 ), .out(\comparator/n46 ) );
  inv \comparator/U45  ( .a(\comparator/N2000 ), .out(\comparator/n45 ) );
  inv \comparator/U44  ( .a(\comparator/N2003 ), .out(\comparator/n44 ) );
  inv \comparator/U43  ( .a(\comparator/N2002 ), .out(\comparator/n43 ) );
  inv \comparator/U42  ( .a(\comparator/N2005 ), .out(\comparator/n42 ) );
  inv \comparator/U41  ( .a(\comparator/N2004 ), .out(\comparator/n41 ) );
  inv \comparator/U40  ( .a(\comparator/N2007 ), .out(\comparator/n40 ) );
  inv \comparator/U39  ( .a(\comparator/N2006 ), .out(\comparator/n39 ) );
  inv \comparator/U38  ( .a(\comparator/N2009 ), .out(\comparator/n38 ) );
  inv \comparator/U37  ( .a(\comparator/N2008 ), .out(\comparator/n37 ) );
  inv \comparator/U36  ( .a(\comparator/N2011 ), .out(\comparator/n36 ) );
  inv \comparator/U35  ( .a(\comparator/N2010 ), .out(\comparator/n35 ) );
  inv \comparator/U34  ( .a(\comparator/N2013 ), .out(\comparator/n34 ) );
  inv \comparator/U33  ( .a(\comparator/N2012 ), .out(\comparator/n33 ) );
  inv \comparator/U32  ( .a(\comparator/N2015 ), .out(\comparator/n32 ) );
  inv \comparator/U31  ( .a(\comparator/N2014 ), .out(\comparator/n31 ) );
  inv \comparator/U30  ( .a(\comparator/N2017 ), .out(\comparator/n30 ) );
  inv \comparator/U29  ( .a(\comparator/N2016 ), .out(\comparator/n29 ) );
  inv \comparator/U28  ( .a(\comparator/N2019 ), .out(\comparator/n28 ) );
  inv \comparator/U27  ( .a(\comparator/N2018 ), .out(\comparator/n27 ) );
  inv \comparator/U26  ( .a(\comparator/N2021 ), .out(\comparator/n26 ) );
  inv \comparator/U25  ( .a(\comparator/N2020 ), .out(\comparator/n25 ) );
  inv \comparator/U24  ( .a(\comparator/N2023 ), .out(\comparator/n24 ) );
  inv \comparator/U23  ( .a(\comparator/N2022 ), .out(\comparator/n23 ) );
  inv \comparator/U22  ( .a(\comparator/N2025 ), .out(\comparator/n22 ) );
  inv \comparator/U21  ( .a(\comparator/N2024 ), .out(\comparator/n21 ) );
  inv \comparator/U20  ( .a(\comparator/N2027 ), .out(\comparator/n20 ) );
  inv \comparator/U19  ( .a(\comparator/N2026 ), .out(\comparator/n19 ) );
  inv \comparator/U18  ( .a(\comparator/N2029 ), .out(\comparator/n18 ) );
  inv \comparator/U17  ( .a(\comparator/N2028 ), .out(\comparator/n17 ) );
  inv \comparator/U16  ( .a(\comparator/N2031 ), .out(\comparator/n16 ) );
  inv \comparator/U15  ( .a(\comparator/N2030 ), .out(\comparator/n15 ) );
  inv \comparator/U14  ( .a(\comparator/N2033 ), .out(\comparator/n14 ) );
  inv \comparator/U13  ( .a(\comparator/N2032 ), .out(\comparator/n13 ) );
  inv \comparator/U12  ( .a(\comparator/N2035 ), .out(\comparator/n12 ) );
  inv \comparator/U11  ( .a(\comparator/N2034 ), .out(\comparator/n11 ) );
  inv \comparator/U10  ( .a(\comparator/N2037 ), .out(\comparator/n10 ) );
  inv \comparator/U9  ( .a(\comparator/N2036 ), .out(\comparator/n9 ) );
  inv \comparator/U8  ( .a(\comparator/N2039 ), .out(\comparator/n8 ) );
  inv \comparator/U7  ( .a(\comparator/N2038 ), .out(\comparator/n7 ) );
  inv \comparator/U6  ( .a(\comparator/N2041 ), .out(\comparator/n6 ) );
  inv \comparator/U5  ( .a(\comparator/N2040 ), .out(\comparator/n5 ) );
  inv \comparator/U4  ( .a(\comparator/N2043 ), .out(\comparator/n4 ) );
  inv \comparator/U3  ( .a(\comparator/N2042 ), .out(\comparator/n3 ) );
  inv \comparator/U2  ( .a(\comparator/N2045 ), .out(\comparator/n2 ) );
  inv \comparator/U1  ( .a(\comparator/N2044 ), .out(\comparator/n1 ) );
  inv \comparator/I_0  ( .a(\comparator/N2046 ), .out(out) );
  nand2 \comparator/C8  ( .a(\comparator/n1 ), .b(\comparator/n2 ), .out(
        \comparator/N2046 ) );
  nand2 \comparator/C9  ( .a(\comparator/n3 ), .b(\comparator/n4 ), .out(
        \comparator/N2044 ) );
  nand2 \comparator/C10  ( .a(\comparator/n5 ), .b(\comparator/n6 ), .out(
        \comparator/N2042 ) );
  nand2 \comparator/C11  ( .a(\comparator/n7 ), .b(\comparator/n8 ), .out(
        \comparator/N2040 ) );
  nand2 \comparator/C12  ( .a(\comparator/n9 ), .b(\comparator/n10 ), .out(
        \comparator/N2038 ) );
  nand2 \comparator/C13  ( .a(\comparator/n11 ), .b(\comparator/n12 ), .out(
        \comparator/N2036 ) );
  nand2 \comparator/C14  ( .a(\comparator/n13 ), .b(\comparator/n14 ), .out(
        \comparator/N2034 ) );
  nand2 \comparator/C15  ( .a(\comparator/n15 ), .b(\comparator/n16 ), .out(
        \comparator/N2032 ) );
  nand2 \comparator/C16  ( .a(\comparator/n17 ), .b(\comparator/n18 ), .out(
        \comparator/N2030 ) );
  nand2 \comparator/C17  ( .a(\comparator/n19 ), .b(\comparator/n20 ), .out(
        \comparator/N2028 ) );
  nand2 \comparator/C18  ( .a(\comparator/n21 ), .b(\comparator/n22 ), .out(
        \comparator/N2026 ) );
  nand2 \comparator/C19  ( .a(\comparator/n23 ), .b(\comparator/n24 ), .out(
        \comparator/N2024 ) );
  nand2 \comparator/C20  ( .a(\comparator/n25 ), .b(\comparator/n26 ), .out(
        \comparator/N2022 ) );
  nand2 \comparator/C21  ( .a(\comparator/n27 ), .b(\comparator/n28 ), .out(
        \comparator/N2020 ) );
  nand2 \comparator/C22  ( .a(\comparator/n29 ), .b(\comparator/n30 ), .out(
        \comparator/N2018 ) );
  nand2 \comparator/C23  ( .a(\comparator/n31 ), .b(\comparator/n32 ), .out(
        \comparator/N2016 ) );
  nand2 \comparator/C24  ( .a(\comparator/n33 ), .b(\comparator/n34 ), .out(
        \comparator/N2014 ) );
  nand2 \comparator/C25  ( .a(\comparator/n35 ), .b(\comparator/n36 ), .out(
        \comparator/N2012 ) );
  nand2 \comparator/C26  ( .a(\comparator/n37 ), .b(\comparator/n38 ), .out(
        \comparator/N2010 ) );
  nand2 \comparator/C27  ( .a(\comparator/n39 ), .b(\comparator/n40 ), .out(
        \comparator/N2008 ) );
  nand2 \comparator/C28  ( .a(\comparator/n41 ), .b(\comparator/n42 ), .out(
        \comparator/N2006 ) );
  nand2 \comparator/C29  ( .a(\comparator/n43 ), .b(\comparator/n44 ), .out(
        \comparator/N2004 ) );
  nand2 \comparator/C30  ( .a(\comparator/n45 ), .b(\comparator/n46 ), .out(
        \comparator/N2002 ) );
  nand2 \comparator/C31  ( .a(\comparator/n47 ), .b(\comparator/n48 ), .out(
        \comparator/N2000 ) );
  nand2 \comparator/C32  ( .a(\comparator/n49 ), .b(\comparator/n50 ), .out(
        \comparator/N1998 ) );
  nand2 \comparator/C33  ( .a(\comparator/n51 ), .b(\comparator/n52 ), .out(
        \comparator/N1996 ) );
  nand2 \comparator/C34  ( .a(\comparator/n53 ), .b(\comparator/n54 ), .out(
        \comparator/N1994 ) );
  nand2 \comparator/C35  ( .a(\comparator/n55 ), .b(\comparator/n56 ), .out(
        \comparator/N1992 ) );
  nand2 \comparator/C36  ( .a(\comparator/n57 ), .b(\comparator/n58 ), .out(
        \comparator/N1990 ) );
  nand2 \comparator/C37  ( .a(\comparator/n59 ), .b(\comparator/n60 ), .out(
        \comparator/N1988 ) );
  nand2 \comparator/C38  ( .a(\comparator/n61 ), .b(\comparator/n62 ), .out(
        \comparator/N1986 ) );
  nand2 \comparator/C39  ( .a(\comparator/n63 ), .b(\comparator/n64 ), .out(
        \comparator/N1984 ) );
  nand2 \comparator/C40  ( .a(\comparator/n65 ), .b(\comparator/n66 ), .out(
        \comparator/N1982 ) );
  nand2 \comparator/C41  ( .a(\comparator/n67 ), .b(\comparator/n68 ), .out(
        \comparator/N1980 ) );
  nand2 \comparator/C42  ( .a(\comparator/n69 ), .b(\comparator/n70 ), .out(
        \comparator/N1978 ) );
  nand2 \comparator/C43  ( .a(\comparator/n71 ), .b(\comparator/n72 ), .out(
        \comparator/N1976 ) );
  nand2 \comparator/C44  ( .a(\comparator/n73 ), .b(\comparator/n74 ), .out(
        \comparator/N1974 ) );
  nand2 \comparator/C45  ( .a(\comparator/n75 ), .b(\comparator/n76 ), .out(
        \comparator/N1972 ) );
  nand2 \comparator/C46  ( .a(\comparator/n77 ), .b(\comparator/n78 ), .out(
        \comparator/N1970 ) );
  nand2 \comparator/C47  ( .a(\comparator/n79 ), .b(\comparator/n80 ), .out(
        \comparator/N1968 ) );
  nand2 \comparator/C48  ( .a(\comparator/n81 ), .b(\comparator/n82 ), .out(
        \comparator/N1966 ) );
  nand2 \comparator/C49  ( .a(\comparator/n83 ), .b(\comparator/n84 ), .out(
        \comparator/N1964 ) );
  nand2 \comparator/C50  ( .a(\comparator/n85 ), .b(\comparator/n86 ), .out(
        \comparator/N1962 ) );
  nand2 \comparator/C51  ( .a(\comparator/n87 ), .b(\comparator/n88 ), .out(
        \comparator/N1960 ) );
  nand2 \comparator/C52  ( .a(\comparator/n89 ), .b(\comparator/n90 ), .out(
        \comparator/N1958 ) );
  nand2 \comparator/C53  ( .a(\comparator/n91 ), .b(\comparator/n92 ), .out(
        \comparator/N1956 ) );
  nand2 \comparator/C54  ( .a(\comparator/n93 ), .b(\comparator/n94 ), .out(
        \comparator/N1954 ) );
  nand2 \comparator/C55  ( .a(\comparator/n95 ), .b(\comparator/n96 ), .out(
        \comparator/N1952 ) );
  nand2 \comparator/C56  ( .a(\comparator/n97 ), .b(\comparator/n98 ), .out(
        \comparator/N1950 ) );
  nand2 \comparator/C57  ( .a(\comparator/n99 ), .b(\comparator/n100 ), .out(
        \comparator/N1948 ) );
  nand2 \comparator/C58  ( .a(\comparator/n101 ), .b(\comparator/n102 ), .out(
        \comparator/N1946 ) );
  nand2 \comparator/C59  ( .a(\comparator/n103 ), .b(\comparator/n104 ), .out(
        \comparator/N1944 ) );
  nand2 \comparator/C60  ( .a(\comparator/n105 ), .b(\comparator/n106 ), .out(
        \comparator/N1942 ) );
  nand2 \comparator/C61  ( .a(\comparator/n107 ), .b(\comparator/n108 ), .out(
        \comparator/N1940 ) );
  nand2 \comparator/C62  ( .a(\comparator/n109 ), .b(\comparator/n110 ), .out(
        \comparator/N1938 ) );
  nand2 \comparator/C63  ( .a(\comparator/n111 ), .b(\comparator/n112 ), .out(
        \comparator/N1936 ) );
  nand2 \comparator/C64  ( .a(\comparator/n113 ), .b(\comparator/n114 ), .out(
        \comparator/N1934 ) );
  nand2 \comparator/C65  ( .a(\comparator/n115 ), .b(\comparator/n116 ), .out(
        \comparator/N1932 ) );
  nand2 \comparator/C66  ( .a(\comparator/n117 ), .b(\comparator/n118 ), .out(
        \comparator/N1930 ) );
  nand2 \comparator/C67  ( .a(\comparator/n119 ), .b(\comparator/n120 ), .out(
        \comparator/N1928 ) );
  nand2 \comparator/C68  ( .a(\comparator/n121 ), .b(\comparator/n122 ), .out(
        \comparator/N1926 ) );
  nand2 \comparator/C69  ( .a(\comparator/n123 ), .b(\comparator/n124 ), .out(
        \comparator/N1924 ) );
  nand2 \comparator/C70  ( .a(\comparator/n125 ), .b(\comparator/n126 ), .out(
        \comparator/N1922 ) );
  nand2 \comparator/C71  ( .a(\comparator/n127 ), .b(\comparator/n128 ), .out(
        \comparator/N1920 ) );
  nand2 \comparator/C72  ( .a(\comparator/n129 ), .b(\comparator/n130 ), .out(
        \comparator/N1918 ) );
  nand2 \comparator/C73  ( .a(\comparator/n131 ), .b(\comparator/n132 ), .out(
        \comparator/N1916 ) );
  nand2 \comparator/C74  ( .a(\comparator/n133 ), .b(\comparator/n134 ), .out(
        \comparator/N1914 ) );
  nand2 \comparator/C75  ( .a(\comparator/n135 ), .b(\comparator/n136 ), .out(
        \comparator/N1912 ) );
  nand2 \comparator/C76  ( .a(\comparator/n137 ), .b(\comparator/n138 ), .out(
        \comparator/N1910 ) );
  nand2 \comparator/C77  ( .a(\comparator/n139 ), .b(\comparator/n140 ), .out(
        \comparator/N1908 ) );
  nand2 \comparator/C78  ( .a(\comparator/n141 ), .b(\comparator/n142 ), .out(
        \comparator/N1906 ) );
  nand2 \comparator/C79  ( .a(\comparator/n143 ), .b(\comparator/n144 ), .out(
        \comparator/N1904 ) );
  nand2 \comparator/C80  ( .a(\comparator/n145 ), .b(\comparator/n146 ), .out(
        \comparator/N1902 ) );
  nand2 \comparator/C81  ( .a(\comparator/n147 ), .b(\comparator/n148 ), .out(
        \comparator/N1900 ) );
  nand2 \comparator/C82  ( .a(\comparator/n149 ), .b(\comparator/n150 ), .out(
        \comparator/N1898 ) );
  nand2 \comparator/C83  ( .a(\comparator/n151 ), .b(\comparator/n152 ), .out(
        \comparator/N1896 ) );
  nand2 \comparator/C84  ( .a(\comparator/n153 ), .b(\comparator/n154 ), .out(
        \comparator/N1894 ) );
  nand2 \comparator/C85  ( .a(\comparator/n155 ), .b(\comparator/n156 ), .out(
        \comparator/N1892 ) );
  nand2 \comparator/C86  ( .a(\comparator/n157 ), .b(\comparator/n158 ), .out(
        \comparator/N1890 ) );
  nand2 \comparator/C87  ( .a(\comparator/n159 ), .b(\comparator/n160 ), .out(
        \comparator/N1888 ) );
  nand2 \comparator/C88  ( .a(\comparator/n161 ), .b(\comparator/n162 ), .out(
        \comparator/N1886 ) );
  nand2 \comparator/C89  ( .a(\comparator/n163 ), .b(\comparator/n164 ), .out(
        \comparator/N1884 ) );
  nand2 \comparator/C90  ( .a(\comparator/n165 ), .b(\comparator/n166 ), .out(
        \comparator/N1882 ) );
  nand2 \comparator/C91  ( .a(\comparator/n167 ), .b(\comparator/n168 ), .out(
        \comparator/N1880 ) );
  nand2 \comparator/C92  ( .a(\comparator/n169 ), .b(\comparator/n170 ), .out(
        \comparator/N1878 ) );
  nand2 \comparator/C93  ( .a(\comparator/n171 ), .b(\comparator/n172 ), .out(
        \comparator/N1876 ) );
  nand2 \comparator/C94  ( .a(\comparator/n173 ), .b(\comparator/n174 ), .out(
        \comparator/N1874 ) );
  nand2 \comparator/C95  ( .a(\comparator/n175 ), .b(\comparator/n176 ), .out(
        \comparator/N1872 ) );
  nand2 \comparator/C96  ( .a(\comparator/n177 ), .b(\comparator/n178 ), .out(
        \comparator/N1870 ) );
  nand2 \comparator/C97  ( .a(\comparator/n179 ), .b(\comparator/n180 ), .out(
        \comparator/N1868 ) );
  nand2 \comparator/C98  ( .a(\comparator/n181 ), .b(\comparator/n182 ), .out(
        \comparator/N1866 ) );
  nand2 \comparator/C99  ( .a(\comparator/n183 ), .b(\comparator/n184 ), .out(
        \comparator/N1864 ) );
  nand2 \comparator/C100  ( .a(\comparator/n185 ), .b(\comparator/n186 ), 
        .out(\comparator/N1862 ) );
  nand2 \comparator/C101  ( .a(\comparator/n187 ), .b(\comparator/n188 ), 
        .out(\comparator/N1860 ) );
  nand2 \comparator/C102  ( .a(\comparator/n189 ), .b(\comparator/n190 ), 
        .out(\comparator/N1858 ) );
  nand2 \comparator/C103  ( .a(\comparator/n191 ), .b(\comparator/n192 ), 
        .out(\comparator/N1856 ) );
  nand2 \comparator/C104  ( .a(\comparator/n193 ), .b(\comparator/n194 ), 
        .out(\comparator/N1854 ) );
  nand2 \comparator/C105  ( .a(\comparator/n195 ), .b(\comparator/n196 ), 
        .out(\comparator/N1852 ) );
  nand2 \comparator/C106  ( .a(\comparator/n197 ), .b(\comparator/n198 ), 
        .out(\comparator/N1850 ) );
  nand2 \comparator/C107  ( .a(\comparator/n199 ), .b(\comparator/n200 ), 
        .out(\comparator/N1848 ) );
  nand2 \comparator/C108  ( .a(\comparator/n201 ), .b(\comparator/n202 ), 
        .out(\comparator/N1846 ) );
  nand2 \comparator/C109  ( .a(\comparator/n203 ), .b(\comparator/n204 ), 
        .out(\comparator/N1844 ) );
  nand2 \comparator/C110  ( .a(\comparator/n205 ), .b(\comparator/n206 ), 
        .out(\comparator/N1842 ) );
  nand2 \comparator/C111  ( .a(\comparator/n207 ), .b(\comparator/n208 ), 
        .out(\comparator/N1840 ) );
  nand2 \comparator/C112  ( .a(\comparator/n209 ), .b(\comparator/n210 ), 
        .out(\comparator/N1838 ) );
  nand2 \comparator/C113  ( .a(\comparator/n211 ), .b(\comparator/n212 ), 
        .out(\comparator/N1836 ) );
  nand2 \comparator/C114  ( .a(\comparator/n213 ), .b(\comparator/n214 ), 
        .out(\comparator/N1834 ) );
  nand2 \comparator/C115  ( .a(\comparator/n215 ), .b(\comparator/n216 ), 
        .out(\comparator/N1832 ) );
  nand2 \comparator/C116  ( .a(\comparator/n217 ), .b(\comparator/n218 ), 
        .out(\comparator/N1830 ) );
  nand2 \comparator/C117  ( .a(\comparator/n219 ), .b(\comparator/n220 ), 
        .out(\comparator/N1828 ) );
  nand2 \comparator/C118  ( .a(\comparator/n221 ), .b(\comparator/n222 ), 
        .out(\comparator/N1826 ) );
  nand2 \comparator/C119  ( .a(\comparator/n223 ), .b(\comparator/n224 ), 
        .out(\comparator/N1824 ) );
  nand2 \comparator/C120  ( .a(\comparator/n225 ), .b(\comparator/n226 ), 
        .out(\comparator/N1822 ) );
  nand2 \comparator/C121  ( .a(\comparator/n227 ), .b(\comparator/n228 ), 
        .out(\comparator/N1820 ) );
  nand2 \comparator/C122  ( .a(\comparator/n229 ), .b(\comparator/n230 ), 
        .out(\comparator/N1818 ) );
  nand2 \comparator/C123  ( .a(\comparator/n231 ), .b(\comparator/n232 ), 
        .out(\comparator/N1816 ) );
  nand2 \comparator/C124  ( .a(\comparator/n233 ), .b(\comparator/n234 ), 
        .out(\comparator/N1814 ) );
  nand2 \comparator/C125  ( .a(\comparator/n235 ), .b(\comparator/n236 ), 
        .out(\comparator/N1812 ) );
  nand2 \comparator/C126  ( .a(\comparator/n237 ), .b(\comparator/n238 ), 
        .out(\comparator/N1810 ) );
  nand2 \comparator/C127  ( .a(\comparator/n239 ), .b(\comparator/n240 ), 
        .out(\comparator/N1808 ) );
  nand2 \comparator/C128  ( .a(\comparator/n241 ), .b(\comparator/n242 ), 
        .out(\comparator/N1806 ) );
  nand2 \comparator/C129  ( .a(\comparator/n243 ), .b(\comparator/n244 ), 
        .out(\comparator/N1804 ) );
  nand2 \comparator/C130  ( .a(\comparator/n245 ), .b(\comparator/n246 ), 
        .out(\comparator/N1802 ) );
  nand2 \comparator/C131  ( .a(\comparator/n247 ), .b(\comparator/n248 ), 
        .out(\comparator/N1800 ) );
  nand2 \comparator/C132  ( .a(\comparator/n249 ), .b(\comparator/n250 ), 
        .out(\comparator/N1798 ) );
  nand2 \comparator/C133  ( .a(\comparator/n251 ), .b(\comparator/n252 ), 
        .out(\comparator/N1796 ) );
  nand2 \comparator/C134  ( .a(\comparator/n253 ), .b(\comparator/n254 ), 
        .out(\comparator/N1794 ) );
  nand2 \comparator/C135  ( .a(\comparator/n255 ), .b(\comparator/n256 ), 
        .out(\comparator/N1792 ) );
  nand2 \comparator/C136  ( .a(\comparator/n257 ), .b(\comparator/n258 ), 
        .out(\comparator/N1790 ) );
  nand2 \comparator/C137  ( .a(\comparator/n259 ), .b(\comparator/n260 ), 
        .out(\comparator/N1788 ) );
  nand2 \comparator/C138  ( .a(\comparator/n261 ), .b(\comparator/n262 ), 
        .out(\comparator/N1786 ) );
  nand2 \comparator/C139  ( .a(\comparator/n263 ), .b(\comparator/n264 ), 
        .out(\comparator/N1784 ) );
  nand2 \comparator/C140  ( .a(\comparator/n265 ), .b(\comparator/n266 ), 
        .out(\comparator/N1782 ) );
  nand2 \comparator/C141  ( .a(\comparator/n267 ), .b(\comparator/n268 ), 
        .out(\comparator/N1780 ) );
  nand2 \comparator/C142  ( .a(\comparator/n269 ), .b(\comparator/n270 ), 
        .out(\comparator/N1778 ) );
  nand2 \comparator/C143  ( .a(\comparator/n271 ), .b(\comparator/n272 ), 
        .out(\comparator/N1776 ) );
  nand2 \comparator/C144  ( .a(\comparator/n273 ), .b(\comparator/n274 ), 
        .out(\comparator/N1774 ) );
  nand2 \comparator/C145  ( .a(\comparator/n275 ), .b(\comparator/n276 ), 
        .out(\comparator/N1772 ) );
  nand2 \comparator/C146  ( .a(\comparator/n277 ), .b(\comparator/n278 ), 
        .out(\comparator/N1770 ) );
  nand2 \comparator/C147  ( .a(\comparator/n279 ), .b(\comparator/n280 ), 
        .out(\comparator/N1768 ) );
  nand2 \comparator/C148  ( .a(\comparator/n281 ), .b(\comparator/n282 ), 
        .out(\comparator/N1766 ) );
  nand2 \comparator/C149  ( .a(\comparator/n283 ), .b(\comparator/n284 ), 
        .out(\comparator/N1764 ) );
  nand2 \comparator/C150  ( .a(\comparator/n285 ), .b(\comparator/n286 ), 
        .out(\comparator/N1762 ) );
  nand2 \comparator/C151  ( .a(\comparator/n287 ), .b(\comparator/n288 ), 
        .out(\comparator/N1760 ) );
  nand2 \comparator/C152  ( .a(\comparator/n289 ), .b(\comparator/n290 ), 
        .out(\comparator/N1758 ) );
  nand2 \comparator/C153  ( .a(\comparator/n291 ), .b(\comparator/n292 ), 
        .out(\comparator/N1756 ) );
  nand2 \comparator/C154  ( .a(\comparator/n293 ), .b(\comparator/n294 ), 
        .out(\comparator/N1754 ) );
  nand2 \comparator/C155  ( .a(\comparator/n295 ), .b(\comparator/n296 ), 
        .out(\comparator/N1752 ) );
  nand2 \comparator/C156  ( .a(\comparator/n297 ), .b(\comparator/n298 ), 
        .out(\comparator/N1750 ) );
  nand2 \comparator/C157  ( .a(\comparator/n299 ), .b(\comparator/n300 ), 
        .out(\comparator/N1748 ) );
  nand2 \comparator/C158  ( .a(\comparator/n301 ), .b(\comparator/n302 ), 
        .out(\comparator/N1746 ) );
  nand2 \comparator/C159  ( .a(\comparator/n303 ), .b(\comparator/n304 ), 
        .out(\comparator/N1744 ) );
  nand2 \comparator/C160  ( .a(\comparator/n305 ), .b(\comparator/n306 ), 
        .out(\comparator/N1742 ) );
  nand2 \comparator/C161  ( .a(\comparator/n307 ), .b(\comparator/n308 ), 
        .out(\comparator/N1740 ) );
  nand2 \comparator/C162  ( .a(\comparator/n309 ), .b(\comparator/n310 ), 
        .out(\comparator/N1738 ) );
  nand2 \comparator/C163  ( .a(\comparator/n311 ), .b(\comparator/n312 ), 
        .out(\comparator/N1736 ) );
  nand2 \comparator/C164  ( .a(\comparator/n313 ), .b(\comparator/n314 ), 
        .out(\comparator/N1734 ) );
  nand2 \comparator/C165  ( .a(\comparator/n315 ), .b(\comparator/n316 ), 
        .out(\comparator/N1732 ) );
  nand2 \comparator/C166  ( .a(\comparator/n317 ), .b(\comparator/n318 ), 
        .out(\comparator/N1730 ) );
  nand2 \comparator/C167  ( .a(\comparator/n319 ), .b(\comparator/n320 ), 
        .out(\comparator/N1728 ) );
  nand2 \comparator/C168  ( .a(\comparator/n321 ), .b(\comparator/n322 ), 
        .out(\comparator/N1726 ) );
  nand2 \comparator/C169  ( .a(\comparator/n323 ), .b(\comparator/n324 ), 
        .out(\comparator/N1724 ) );
  nand2 \comparator/C170  ( .a(\comparator/n325 ), .b(\comparator/n326 ), 
        .out(\comparator/N1722 ) );
  nand2 \comparator/C171  ( .a(\comparator/n327 ), .b(\comparator/n328 ), 
        .out(\comparator/N1720 ) );
  nand2 \comparator/C172  ( .a(\comparator/n329 ), .b(\comparator/n330 ), 
        .out(\comparator/N1718 ) );
  nand2 \comparator/C173  ( .a(\comparator/n331 ), .b(\comparator/n332 ), 
        .out(\comparator/N1716 ) );
  nand2 \comparator/C174  ( .a(\comparator/n333 ), .b(\comparator/n334 ), 
        .out(\comparator/N1714 ) );
  nand2 \comparator/C175  ( .a(\comparator/n335 ), .b(\comparator/n336 ), 
        .out(\comparator/N1712 ) );
  nand2 \comparator/C176  ( .a(\comparator/n337 ), .b(\comparator/n338 ), 
        .out(\comparator/N1710 ) );
  nand2 \comparator/C177  ( .a(\comparator/n339 ), .b(\comparator/n340 ), 
        .out(\comparator/N1708 ) );
  nand2 \comparator/C178  ( .a(\comparator/n341 ), .b(\comparator/n342 ), 
        .out(\comparator/N1706 ) );
  nand2 \comparator/C179  ( .a(\comparator/n343 ), .b(\comparator/n344 ), 
        .out(\comparator/N1704 ) );
  nand2 \comparator/C180  ( .a(\comparator/n345 ), .b(\comparator/n346 ), 
        .out(\comparator/N1702 ) );
  nand2 \comparator/C181  ( .a(\comparator/n347 ), .b(\comparator/n348 ), 
        .out(\comparator/N1700 ) );
  nand2 \comparator/C182  ( .a(\comparator/n349 ), .b(\comparator/n350 ), 
        .out(\comparator/N1698 ) );
  nand2 \comparator/C183  ( .a(\comparator/n351 ), .b(\comparator/n352 ), 
        .out(\comparator/N1696 ) );
  nand2 \comparator/C184  ( .a(\comparator/n353 ), .b(\comparator/n354 ), 
        .out(\comparator/N1694 ) );
  nand2 \comparator/C185  ( .a(\comparator/n355 ), .b(\comparator/n356 ), 
        .out(\comparator/N1692 ) );
  nand2 \comparator/C186  ( .a(\comparator/n357 ), .b(\comparator/n358 ), 
        .out(\comparator/N1690 ) );
  nand2 \comparator/C187  ( .a(\comparator/n359 ), .b(\comparator/n360 ), 
        .out(\comparator/N1688 ) );
  nand2 \comparator/C188  ( .a(\comparator/n361 ), .b(\comparator/n362 ), 
        .out(\comparator/N1686 ) );
  nand2 \comparator/C189  ( .a(\comparator/n363 ), .b(\comparator/n364 ), 
        .out(\comparator/N1684 ) );
  nand2 \comparator/C190  ( .a(\comparator/n365 ), .b(\comparator/n366 ), 
        .out(\comparator/N1682 ) );
  nand2 \comparator/C191  ( .a(\comparator/n367 ), .b(\comparator/n368 ), 
        .out(\comparator/N1680 ) );
  nand2 \comparator/C192  ( .a(\comparator/n369 ), .b(\comparator/n370 ), 
        .out(\comparator/N1678 ) );
  nand2 \comparator/C193  ( .a(\comparator/n371 ), .b(\comparator/n372 ), 
        .out(\comparator/N1676 ) );
  nand2 \comparator/C194  ( .a(\comparator/n373 ), .b(\comparator/n374 ), 
        .out(\comparator/N1674 ) );
  nand2 \comparator/C195  ( .a(\comparator/n375 ), .b(\comparator/n376 ), 
        .out(\comparator/N1672 ) );
  nand2 \comparator/C196  ( .a(\comparator/n377 ), .b(\comparator/n378 ), 
        .out(\comparator/N1670 ) );
  nand2 \comparator/C197  ( .a(\comparator/n379 ), .b(\comparator/n380 ), 
        .out(\comparator/N1668 ) );
  nand2 \comparator/C198  ( .a(\comparator/n381 ), .b(\comparator/n382 ), 
        .out(\comparator/N1666 ) );
  nand2 \comparator/C199  ( .a(\comparator/n383 ), .b(\comparator/n384 ), 
        .out(\comparator/N1664 ) );
  nand2 \comparator/C200  ( .a(\comparator/n385 ), .b(\comparator/n386 ), 
        .out(\comparator/N1662 ) );
  nand2 \comparator/C201  ( .a(\comparator/n387 ), .b(\comparator/n388 ), 
        .out(\comparator/N1660 ) );
  nand2 \comparator/C202  ( .a(\comparator/n389 ), .b(\comparator/n390 ), 
        .out(\comparator/N1658 ) );
  nand2 \comparator/C203  ( .a(\comparator/n391 ), .b(\comparator/n392 ), 
        .out(\comparator/N1656 ) );
  nand2 \comparator/C204  ( .a(\comparator/n393 ), .b(\comparator/n394 ), 
        .out(\comparator/N1654 ) );
  nand2 \comparator/C205  ( .a(\comparator/n395 ), .b(\comparator/n396 ), 
        .out(\comparator/N1652 ) );
  nand2 \comparator/C206  ( .a(\comparator/n397 ), .b(\comparator/n398 ), 
        .out(\comparator/N1650 ) );
  nand2 \comparator/C207  ( .a(\comparator/n399 ), .b(\comparator/n400 ), 
        .out(\comparator/N1648 ) );
  nand2 \comparator/C208  ( .a(\comparator/n401 ), .b(\comparator/n402 ), 
        .out(\comparator/N1646 ) );
  nand2 \comparator/C209  ( .a(\comparator/n403 ), .b(\comparator/n404 ), 
        .out(\comparator/N1644 ) );
  nand2 \comparator/C210  ( .a(\comparator/n405 ), .b(\comparator/n406 ), 
        .out(\comparator/N1642 ) );
  nand2 \comparator/C211  ( .a(\comparator/n407 ), .b(\comparator/n408 ), 
        .out(\comparator/N1640 ) );
  nand2 \comparator/C212  ( .a(\comparator/n409 ), .b(\comparator/n410 ), 
        .out(\comparator/N1638 ) );
  nand2 \comparator/C213  ( .a(\comparator/n411 ), .b(\comparator/n412 ), 
        .out(\comparator/N1636 ) );
  nand2 \comparator/C214  ( .a(\comparator/n413 ), .b(\comparator/n414 ), 
        .out(\comparator/N1634 ) );
  nand2 \comparator/C215  ( .a(\comparator/n415 ), .b(\comparator/n416 ), 
        .out(\comparator/N1632 ) );
  nand2 \comparator/C216  ( .a(\comparator/n417 ), .b(\comparator/n418 ), 
        .out(\comparator/N1630 ) );
  nand2 \comparator/C217  ( .a(\comparator/n419 ), .b(\comparator/n420 ), 
        .out(\comparator/N1628 ) );
  nand2 \comparator/C218  ( .a(\comparator/n421 ), .b(\comparator/n422 ), 
        .out(\comparator/N1626 ) );
  nand2 \comparator/C219  ( .a(\comparator/n423 ), .b(\comparator/n424 ), 
        .out(\comparator/N1624 ) );
  nand2 \comparator/C220  ( .a(\comparator/n425 ), .b(\comparator/n426 ), 
        .out(\comparator/N1622 ) );
  nand2 \comparator/C221  ( .a(\comparator/n427 ), .b(\comparator/n428 ), 
        .out(\comparator/N1620 ) );
  nand2 \comparator/C222  ( .a(\comparator/n429 ), .b(\comparator/n430 ), 
        .out(\comparator/N1618 ) );
  nand2 \comparator/C223  ( .a(\comparator/n431 ), .b(\comparator/n432 ), 
        .out(\comparator/N1616 ) );
  nand2 \comparator/C224  ( .a(\comparator/n433 ), .b(\comparator/n434 ), 
        .out(\comparator/N1614 ) );
  nand2 \comparator/C225  ( .a(\comparator/n435 ), .b(\comparator/n436 ), 
        .out(\comparator/N1612 ) );
  nand2 \comparator/C226  ( .a(\comparator/n437 ), .b(\comparator/n438 ), 
        .out(\comparator/N1610 ) );
  nand2 \comparator/C227  ( .a(\comparator/n439 ), .b(\comparator/n440 ), 
        .out(\comparator/N1608 ) );
  nand2 \comparator/C228  ( .a(\comparator/n441 ), .b(\comparator/n442 ), 
        .out(\comparator/N1606 ) );
  nand2 \comparator/C229  ( .a(\comparator/n443 ), .b(\comparator/n444 ), 
        .out(\comparator/N1604 ) );
  nand2 \comparator/C230  ( .a(\comparator/n445 ), .b(\comparator/n446 ), 
        .out(\comparator/N1602 ) );
  nand2 \comparator/C231  ( .a(\comparator/n447 ), .b(\comparator/n448 ), 
        .out(\comparator/N1600 ) );
  nand2 \comparator/C232  ( .a(\comparator/n449 ), .b(\comparator/n450 ), 
        .out(\comparator/N1598 ) );
  nand2 \comparator/C233  ( .a(\comparator/n451 ), .b(\comparator/n452 ), 
        .out(\comparator/N1596 ) );
  nand2 \comparator/C234  ( .a(\comparator/n453 ), .b(\comparator/n454 ), 
        .out(\comparator/N1594 ) );
  nand2 \comparator/C235  ( .a(\comparator/n455 ), .b(\comparator/n456 ), 
        .out(\comparator/N1592 ) );
  nand2 \comparator/C236  ( .a(\comparator/n457 ), .b(\comparator/n458 ), 
        .out(\comparator/N1590 ) );
  nand2 \comparator/C237  ( .a(\comparator/n459 ), .b(\comparator/n460 ), 
        .out(\comparator/N1588 ) );
  nand2 \comparator/C238  ( .a(\comparator/n461 ), .b(\comparator/n462 ), 
        .out(\comparator/N1586 ) );
  nand2 \comparator/C239  ( .a(\comparator/n463 ), .b(\comparator/n464 ), 
        .out(\comparator/N1584 ) );
  nand2 \comparator/C240  ( .a(\comparator/n465 ), .b(\comparator/n466 ), 
        .out(\comparator/N1582 ) );
  nand2 \comparator/C241  ( .a(\comparator/n467 ), .b(\comparator/n468 ), 
        .out(\comparator/N1580 ) );
  nand2 \comparator/C242  ( .a(\comparator/n469 ), .b(\comparator/n470 ), 
        .out(\comparator/N1578 ) );
  nand2 \comparator/C243  ( .a(\comparator/n471 ), .b(\comparator/n472 ), 
        .out(\comparator/N1576 ) );
  nand2 \comparator/C244  ( .a(\comparator/n473 ), .b(\comparator/n474 ), 
        .out(\comparator/N1574 ) );
  nand2 \comparator/C245  ( .a(\comparator/n475 ), .b(\comparator/n476 ), 
        .out(\comparator/N1572 ) );
  nand2 \comparator/C246  ( .a(\comparator/n477 ), .b(\comparator/n478 ), 
        .out(\comparator/N1570 ) );
  nand2 \comparator/C247  ( .a(\comparator/n479 ), .b(\comparator/n480 ), 
        .out(\comparator/N1568 ) );
  nand2 \comparator/C248  ( .a(\comparator/n481 ), .b(\comparator/n482 ), 
        .out(\comparator/N1566 ) );
  nand2 \comparator/C249  ( .a(\comparator/n483 ), .b(\comparator/n484 ), 
        .out(\comparator/N1564 ) );
  nand2 \comparator/C250  ( .a(\comparator/n485 ), .b(\comparator/n486 ), 
        .out(\comparator/N1562 ) );
  nand2 \comparator/C251  ( .a(\comparator/n487 ), .b(\comparator/n488 ), 
        .out(\comparator/N1560 ) );
  nand2 \comparator/C252  ( .a(\comparator/n489 ), .b(\comparator/n490 ), 
        .out(\comparator/N1558 ) );
  nand2 \comparator/C253  ( .a(\comparator/n491 ), .b(\comparator/n492 ), 
        .out(\comparator/N1556 ) );
  nand2 \comparator/C254  ( .a(\comparator/n493 ), .b(\comparator/n494 ), 
        .out(\comparator/N1554 ) );
  nand2 \comparator/C255  ( .a(\comparator/n495 ), .b(\comparator/n496 ), 
        .out(\comparator/N1552 ) );
  nand2 \comparator/C256  ( .a(\comparator/n497 ), .b(\comparator/n498 ), 
        .out(\comparator/N1550 ) );
  nand2 \comparator/C257  ( .a(\comparator/n499 ), .b(\comparator/n500 ), 
        .out(\comparator/N1548 ) );
  nand2 \comparator/C258  ( .a(\comparator/n501 ), .b(\comparator/n502 ), 
        .out(\comparator/N1546 ) );
  nand2 \comparator/C259  ( .a(\comparator/n503 ), .b(\comparator/n504 ), 
        .out(\comparator/N1544 ) );
  nand2 \comparator/C260  ( .a(\comparator/n505 ), .b(\comparator/n506 ), 
        .out(\comparator/N1542 ) );
  nand2 \comparator/C261  ( .a(\comparator/n507 ), .b(\comparator/n508 ), 
        .out(\comparator/N1540 ) );
  nand2 \comparator/C262  ( .a(\comparator/n509 ), .b(\comparator/n510 ), 
        .out(\comparator/N1538 ) );
  nand2 \comparator/C263  ( .a(\comparator/n511 ), .b(\comparator/n512 ), 
        .out(\comparator/N1536 ) );
  nand2 \comparator/C264  ( .a(\comparator/n513 ), .b(\comparator/n514 ), 
        .out(\comparator/N1534 ) );
  nand2 \comparator/C265  ( .a(\comparator/n515 ), .b(\comparator/n516 ), 
        .out(\comparator/N1532 ) );
  nand2 \comparator/C266  ( .a(\comparator/n517 ), .b(\comparator/n518 ), 
        .out(\comparator/N1530 ) );
  nand2 \comparator/C267  ( .a(\comparator/n519 ), .b(\comparator/n520 ), 
        .out(\comparator/N1528 ) );
  nand2 \comparator/C268  ( .a(\comparator/n521 ), .b(\comparator/n522 ), 
        .out(\comparator/N1526 ) );
  nand2 \comparator/C269  ( .a(\comparator/n523 ), .b(\comparator/n524 ), 
        .out(\comparator/N1524 ) );
  nand2 \comparator/C270  ( .a(\comparator/n525 ), .b(\comparator/n526 ), 
        .out(\comparator/N1522 ) );
  nand2 \comparator/C271  ( .a(\comparator/n527 ), .b(\comparator/n528 ), 
        .out(\comparator/N1520 ) );
  nand2 \comparator/C272  ( .a(\comparator/n529 ), .b(\comparator/n530 ), 
        .out(\comparator/N1518 ) );
  nand2 \comparator/C273  ( .a(\comparator/n531 ), .b(\comparator/n532 ), 
        .out(\comparator/N1516 ) );
  nand2 \comparator/C274  ( .a(\comparator/n533 ), .b(\comparator/n534 ), 
        .out(\comparator/N1514 ) );
  nand2 \comparator/C275  ( .a(\comparator/n535 ), .b(\comparator/n536 ), 
        .out(\comparator/N1512 ) );
  nand2 \comparator/C276  ( .a(\comparator/n537 ), .b(\comparator/n538 ), 
        .out(\comparator/N1510 ) );
  nand2 \comparator/C277  ( .a(\comparator/n539 ), .b(\comparator/n540 ), 
        .out(\comparator/N1508 ) );
  nand2 \comparator/C278  ( .a(\comparator/n541 ), .b(\comparator/n542 ), 
        .out(\comparator/N1506 ) );
  nand2 \comparator/C279  ( .a(\comparator/n543 ), .b(\comparator/n544 ), 
        .out(\comparator/N1504 ) );
  nand2 \comparator/C280  ( .a(\comparator/n545 ), .b(\comparator/n546 ), 
        .out(\comparator/N1502 ) );
  nand2 \comparator/C281  ( .a(\comparator/n547 ), .b(\comparator/n548 ), 
        .out(\comparator/N1500 ) );
  nand2 \comparator/C282  ( .a(\comparator/n549 ), .b(\comparator/n550 ), 
        .out(\comparator/N1498 ) );
  nand2 \comparator/C283  ( .a(\comparator/n551 ), .b(\comparator/n552 ), 
        .out(\comparator/N1496 ) );
  nand2 \comparator/C284  ( .a(\comparator/n553 ), .b(\comparator/n554 ), 
        .out(\comparator/N1494 ) );
  nand2 \comparator/C285  ( .a(\comparator/n555 ), .b(\comparator/n556 ), 
        .out(\comparator/N1492 ) );
  nand2 \comparator/C286  ( .a(\comparator/n557 ), .b(\comparator/n558 ), 
        .out(\comparator/N1490 ) );
  nand2 \comparator/C287  ( .a(\comparator/n559 ), .b(\comparator/n560 ), 
        .out(\comparator/N1488 ) );
  nand2 \comparator/C288  ( .a(\comparator/n561 ), .b(\comparator/n562 ), 
        .out(\comparator/N1486 ) );
  nand2 \comparator/C289  ( .a(\comparator/n563 ), .b(\comparator/n564 ), 
        .out(\comparator/N1484 ) );
  nand2 \comparator/C290  ( .a(\comparator/n565 ), .b(\comparator/n566 ), 
        .out(\comparator/N1482 ) );
  nand2 \comparator/C291  ( .a(\comparator/n567 ), .b(\comparator/n568 ), 
        .out(\comparator/N1480 ) );
  nand2 \comparator/C292  ( .a(\comparator/n569 ), .b(\comparator/n570 ), 
        .out(\comparator/N1478 ) );
  nand2 \comparator/C293  ( .a(\comparator/n571 ), .b(\comparator/n572 ), 
        .out(\comparator/N1476 ) );
  nand2 \comparator/C294  ( .a(\comparator/n573 ), .b(\comparator/n574 ), 
        .out(\comparator/N1474 ) );
  nand2 \comparator/C295  ( .a(\comparator/n575 ), .b(\comparator/n576 ), 
        .out(\comparator/N1472 ) );
  nand2 \comparator/C296  ( .a(\comparator/n577 ), .b(\comparator/n578 ), 
        .out(\comparator/N1470 ) );
  nand2 \comparator/C297  ( .a(\comparator/n579 ), .b(\comparator/n580 ), 
        .out(\comparator/N1468 ) );
  nand2 \comparator/C298  ( .a(\comparator/n581 ), .b(\comparator/n582 ), 
        .out(\comparator/N1466 ) );
  nand2 \comparator/C299  ( .a(\comparator/n583 ), .b(\comparator/n584 ), 
        .out(\comparator/N1464 ) );
  nand2 \comparator/C300  ( .a(\comparator/n585 ), .b(\comparator/n586 ), 
        .out(\comparator/N1462 ) );
  nand2 \comparator/C301  ( .a(\comparator/n587 ), .b(\comparator/n588 ), 
        .out(\comparator/N1460 ) );
  nand2 \comparator/C302  ( .a(\comparator/n589 ), .b(\comparator/n590 ), 
        .out(\comparator/N1458 ) );
  nand2 \comparator/C303  ( .a(\comparator/n591 ), .b(\comparator/n592 ), 
        .out(\comparator/N1456 ) );
  nand2 \comparator/C304  ( .a(\comparator/n593 ), .b(\comparator/n594 ), 
        .out(\comparator/N1454 ) );
  nand2 \comparator/C305  ( .a(\comparator/n595 ), .b(\comparator/n596 ), 
        .out(\comparator/N1452 ) );
  nand2 \comparator/C306  ( .a(\comparator/n597 ), .b(\comparator/n598 ), 
        .out(\comparator/N1450 ) );
  nand2 \comparator/C307  ( .a(\comparator/n599 ), .b(\comparator/n600 ), 
        .out(\comparator/N1448 ) );
  nand2 \comparator/C308  ( .a(\comparator/n601 ), .b(\comparator/n602 ), 
        .out(\comparator/N1446 ) );
  nand2 \comparator/C309  ( .a(\comparator/n603 ), .b(\comparator/n604 ), 
        .out(\comparator/N1444 ) );
  nand2 \comparator/C310  ( .a(\comparator/n605 ), .b(\comparator/n606 ), 
        .out(\comparator/N1442 ) );
  nand2 \comparator/C311  ( .a(\comparator/n607 ), .b(\comparator/n608 ), 
        .out(\comparator/N1440 ) );
  nand2 \comparator/C312  ( .a(\comparator/n609 ), .b(\comparator/n610 ), 
        .out(\comparator/N1438 ) );
  nand2 \comparator/C313  ( .a(\comparator/n611 ), .b(\comparator/n612 ), 
        .out(\comparator/N1436 ) );
  nand2 \comparator/C314  ( .a(\comparator/n613 ), .b(\comparator/n614 ), 
        .out(\comparator/N1434 ) );
  nand2 \comparator/C315  ( .a(\comparator/n615 ), .b(\comparator/n616 ), 
        .out(\comparator/N1432 ) );
  nand2 \comparator/C316  ( .a(\comparator/n617 ), .b(\comparator/n618 ), 
        .out(\comparator/N1430 ) );
  nand2 \comparator/C317  ( .a(\comparator/n619 ), .b(\comparator/n620 ), 
        .out(\comparator/N1428 ) );
  nand2 \comparator/C318  ( .a(\comparator/n621 ), .b(\comparator/n622 ), 
        .out(\comparator/N1426 ) );
  nand2 \comparator/C319  ( .a(\comparator/n623 ), .b(\comparator/n624 ), 
        .out(\comparator/N1424 ) );
  nand2 \comparator/C320  ( .a(\comparator/n625 ), .b(\comparator/n626 ), 
        .out(\comparator/N1422 ) );
  nand2 \comparator/C321  ( .a(\comparator/n627 ), .b(\comparator/n628 ), 
        .out(\comparator/N1420 ) );
  nand2 \comparator/C322  ( .a(\comparator/n629 ), .b(\comparator/n630 ), 
        .out(\comparator/N1418 ) );
  nand2 \comparator/C323  ( .a(\comparator/n631 ), .b(\comparator/n632 ), 
        .out(\comparator/N1416 ) );
  nand2 \comparator/C324  ( .a(\comparator/n633 ), .b(\comparator/n634 ), 
        .out(\comparator/N1414 ) );
  nand2 \comparator/C325  ( .a(\comparator/n635 ), .b(\comparator/n636 ), 
        .out(\comparator/N1412 ) );
  nand2 \comparator/C326  ( .a(\comparator/n637 ), .b(\comparator/n638 ), 
        .out(\comparator/N1410 ) );
  nand2 \comparator/C327  ( .a(\comparator/n639 ), .b(\comparator/n640 ), 
        .out(\comparator/N1408 ) );
  nand2 \comparator/C328  ( .a(\comparator/n641 ), .b(\comparator/n642 ), 
        .out(\comparator/N1406 ) );
  nand2 \comparator/C329  ( .a(\comparator/n643 ), .b(\comparator/n644 ), 
        .out(\comparator/N1404 ) );
  nand2 \comparator/C330  ( .a(\comparator/n645 ), .b(\comparator/n646 ), 
        .out(\comparator/N1402 ) );
  nand2 \comparator/C331  ( .a(\comparator/n647 ), .b(\comparator/n648 ), 
        .out(\comparator/N1400 ) );
  nand2 \comparator/C332  ( .a(\comparator/n649 ), .b(\comparator/n650 ), 
        .out(\comparator/N1398 ) );
  nand2 \comparator/C333  ( .a(\comparator/n651 ), .b(\comparator/n652 ), 
        .out(\comparator/N1396 ) );
  nand2 \comparator/C334  ( .a(\comparator/n653 ), .b(\comparator/n654 ), 
        .out(\comparator/N1394 ) );
  nand2 \comparator/C335  ( .a(\comparator/n655 ), .b(\comparator/n656 ), 
        .out(\comparator/N1392 ) );
  nand2 \comparator/C336  ( .a(\comparator/n657 ), .b(\comparator/n658 ), 
        .out(\comparator/N1390 ) );
  nand2 \comparator/C337  ( .a(\comparator/n659 ), .b(\comparator/n660 ), 
        .out(\comparator/N1388 ) );
  nand2 \comparator/C338  ( .a(\comparator/n661 ), .b(\comparator/n662 ), 
        .out(\comparator/N1386 ) );
  nand2 \comparator/C339  ( .a(\comparator/n663 ), .b(\comparator/n664 ), 
        .out(\comparator/N1384 ) );
  nand2 \comparator/C340  ( .a(\comparator/n665 ), .b(\comparator/n666 ), 
        .out(\comparator/N1382 ) );
  nand2 \comparator/C341  ( .a(\comparator/n667 ), .b(\comparator/n668 ), 
        .out(\comparator/N1380 ) );
  nand2 \comparator/C342  ( .a(\comparator/n669 ), .b(\comparator/n670 ), 
        .out(\comparator/N1378 ) );
  nand2 \comparator/C343  ( .a(\comparator/n671 ), .b(\comparator/n672 ), 
        .out(\comparator/N1376 ) );
  nand2 \comparator/C344  ( .a(\comparator/n673 ), .b(\comparator/n674 ), 
        .out(\comparator/N1374 ) );
  nand2 \comparator/C345  ( .a(\comparator/n675 ), .b(\comparator/n676 ), 
        .out(\comparator/N1372 ) );
  nand2 \comparator/C346  ( .a(\comparator/n677 ), .b(\comparator/n678 ), 
        .out(\comparator/N1370 ) );
  nand2 \comparator/C347  ( .a(\comparator/n679 ), .b(\comparator/n680 ), 
        .out(\comparator/N1368 ) );
  nand2 \comparator/C348  ( .a(\comparator/n681 ), .b(\comparator/n682 ), 
        .out(\comparator/N1366 ) );
  nand2 \comparator/C349  ( .a(\comparator/n683 ), .b(\comparator/n684 ), 
        .out(\comparator/N1364 ) );
  nand2 \comparator/C350  ( .a(\comparator/n685 ), .b(\comparator/n686 ), 
        .out(\comparator/N1362 ) );
  nand2 \comparator/C351  ( .a(\comparator/n687 ), .b(\comparator/n688 ), 
        .out(\comparator/N1360 ) );
  nand2 \comparator/C352  ( .a(\comparator/n689 ), .b(\comparator/n690 ), 
        .out(\comparator/N1358 ) );
  nand2 \comparator/C353  ( .a(\comparator/n691 ), .b(\comparator/n692 ), 
        .out(\comparator/N1356 ) );
  nand2 \comparator/C354  ( .a(\comparator/n693 ), .b(\comparator/n694 ), 
        .out(\comparator/N1354 ) );
  nand2 \comparator/C355  ( .a(\comparator/n695 ), .b(\comparator/n696 ), 
        .out(\comparator/N1352 ) );
  nand2 \comparator/C356  ( .a(\comparator/n697 ), .b(\comparator/n698 ), 
        .out(\comparator/N1350 ) );
  nand2 \comparator/C357  ( .a(\comparator/n699 ), .b(\comparator/n700 ), 
        .out(\comparator/N1348 ) );
  nand2 \comparator/C358  ( .a(\comparator/n701 ), .b(\comparator/n702 ), 
        .out(\comparator/N1346 ) );
  nand2 \comparator/C359  ( .a(\comparator/n703 ), .b(\comparator/n704 ), 
        .out(\comparator/N1344 ) );
  nand2 \comparator/C360  ( .a(\comparator/n705 ), .b(\comparator/n706 ), 
        .out(\comparator/N1342 ) );
  nand2 \comparator/C361  ( .a(\comparator/n707 ), .b(\comparator/n708 ), 
        .out(\comparator/N1340 ) );
  nand2 \comparator/C362  ( .a(\comparator/n709 ), .b(\comparator/n710 ), 
        .out(\comparator/N1338 ) );
  nand2 \comparator/C363  ( .a(\comparator/n711 ), .b(\comparator/n712 ), 
        .out(\comparator/N1336 ) );
  nand2 \comparator/C364  ( .a(\comparator/n713 ), .b(\comparator/n714 ), 
        .out(\comparator/N1334 ) );
  nand2 \comparator/C365  ( .a(\comparator/n715 ), .b(\comparator/n716 ), 
        .out(\comparator/N1332 ) );
  nand2 \comparator/C366  ( .a(\comparator/n717 ), .b(\comparator/n718 ), 
        .out(\comparator/N1330 ) );
  nand2 \comparator/C367  ( .a(\comparator/n719 ), .b(\comparator/n720 ), 
        .out(\comparator/N1328 ) );
  nand2 \comparator/C368  ( .a(\comparator/n721 ), .b(\comparator/n722 ), 
        .out(\comparator/N1326 ) );
  nand2 \comparator/C369  ( .a(\comparator/n723 ), .b(\comparator/n724 ), 
        .out(\comparator/N1324 ) );
  nand2 \comparator/C370  ( .a(\comparator/n725 ), .b(\comparator/n726 ), 
        .out(\comparator/N1322 ) );
  nand2 \comparator/C371  ( .a(\comparator/n727 ), .b(\comparator/n728 ), 
        .out(\comparator/N1320 ) );
  nand2 \comparator/C372  ( .a(\comparator/n729 ), .b(\comparator/n730 ), 
        .out(\comparator/N1318 ) );
  nand2 \comparator/C373  ( .a(\comparator/n731 ), .b(\comparator/n732 ), 
        .out(\comparator/N1316 ) );
  nand2 \comparator/C374  ( .a(\comparator/n733 ), .b(\comparator/n734 ), 
        .out(\comparator/N1314 ) );
  nand2 \comparator/C375  ( .a(\comparator/n735 ), .b(\comparator/n736 ), 
        .out(\comparator/N1312 ) );
  nand2 \comparator/C376  ( .a(\comparator/n737 ), .b(\comparator/n738 ), 
        .out(\comparator/N1310 ) );
  nand2 \comparator/C377  ( .a(\comparator/n739 ), .b(\comparator/n740 ), 
        .out(\comparator/N1308 ) );
  nand2 \comparator/C378  ( .a(\comparator/n741 ), .b(\comparator/n742 ), 
        .out(\comparator/N1306 ) );
  nand2 \comparator/C379  ( .a(\comparator/n743 ), .b(\comparator/n744 ), 
        .out(\comparator/N1304 ) );
  nand2 \comparator/C380  ( .a(\comparator/n745 ), .b(\comparator/n746 ), 
        .out(\comparator/N1302 ) );
  nand2 \comparator/C381  ( .a(\comparator/n747 ), .b(\comparator/n748 ), 
        .out(\comparator/N1300 ) );
  nand2 \comparator/C382  ( .a(\comparator/n749 ), .b(\comparator/n750 ), 
        .out(\comparator/N1298 ) );
  nand2 \comparator/C383  ( .a(\comparator/n751 ), .b(\comparator/n752 ), 
        .out(\comparator/N1296 ) );
  nand2 \comparator/C384  ( .a(\comparator/n753 ), .b(\comparator/n754 ), 
        .out(\comparator/N1294 ) );
  nand2 \comparator/C385  ( .a(\comparator/n755 ), .b(\comparator/n756 ), 
        .out(\comparator/N1292 ) );
  nand2 \comparator/C386  ( .a(\comparator/n757 ), .b(\comparator/n758 ), 
        .out(\comparator/N1290 ) );
  nand2 \comparator/C387  ( .a(\comparator/n759 ), .b(\comparator/n760 ), 
        .out(\comparator/N1288 ) );
  nand2 \comparator/C388  ( .a(\comparator/n761 ), .b(\comparator/n762 ), 
        .out(\comparator/N1286 ) );
  nand2 \comparator/C389  ( .a(\comparator/n763 ), .b(\comparator/n764 ), 
        .out(\comparator/N1284 ) );
  nand2 \comparator/C390  ( .a(\comparator/n765 ), .b(\comparator/n766 ), 
        .out(\comparator/N1282 ) );
  nand2 \comparator/C391  ( .a(\comparator/n767 ), .b(\comparator/n768 ), 
        .out(\comparator/N1280 ) );
  nand2 \comparator/C392  ( .a(\comparator/n769 ), .b(\comparator/n770 ), 
        .out(\comparator/N1278 ) );
  nand2 \comparator/C393  ( .a(\comparator/n771 ), .b(\comparator/n772 ), 
        .out(\comparator/N1276 ) );
  nand2 \comparator/C394  ( .a(\comparator/n773 ), .b(\comparator/n774 ), 
        .out(\comparator/N1274 ) );
  nand2 \comparator/C395  ( .a(\comparator/n775 ), .b(\comparator/n776 ), 
        .out(\comparator/N1272 ) );
  nand2 \comparator/C396  ( .a(\comparator/n777 ), .b(\comparator/n778 ), 
        .out(\comparator/N1270 ) );
  nand2 \comparator/C397  ( .a(\comparator/n779 ), .b(\comparator/n780 ), 
        .out(\comparator/N1268 ) );
  nand2 \comparator/C398  ( .a(\comparator/n781 ), .b(\comparator/n782 ), 
        .out(\comparator/N1266 ) );
  nand2 \comparator/C399  ( .a(\comparator/n783 ), .b(\comparator/n784 ), 
        .out(\comparator/N1264 ) );
  nand2 \comparator/C400  ( .a(\comparator/n785 ), .b(\comparator/n786 ), 
        .out(\comparator/N1262 ) );
  nand2 \comparator/C401  ( .a(\comparator/n787 ), .b(\comparator/n788 ), 
        .out(\comparator/N1260 ) );
  nand2 \comparator/C402  ( .a(\comparator/n789 ), .b(\comparator/n790 ), 
        .out(\comparator/N1258 ) );
  nand2 \comparator/C403  ( .a(\comparator/n791 ), .b(\comparator/n792 ), 
        .out(\comparator/N1256 ) );
  nand2 \comparator/C404  ( .a(\comparator/n793 ), .b(\comparator/n794 ), 
        .out(\comparator/N1254 ) );
  nand2 \comparator/C405  ( .a(\comparator/n795 ), .b(\comparator/n796 ), 
        .out(\comparator/N1252 ) );
  nand2 \comparator/C406  ( .a(\comparator/n797 ), .b(\comparator/n798 ), 
        .out(\comparator/N1250 ) );
  nand2 \comparator/C407  ( .a(\comparator/n799 ), .b(\comparator/n800 ), 
        .out(\comparator/N1248 ) );
  nand2 \comparator/C408  ( .a(\comparator/n801 ), .b(\comparator/n802 ), 
        .out(\comparator/N1246 ) );
  nand2 \comparator/C409  ( .a(\comparator/n803 ), .b(\comparator/n804 ), 
        .out(\comparator/N1244 ) );
  nand2 \comparator/C410  ( .a(\comparator/n805 ), .b(\comparator/n806 ), 
        .out(\comparator/N1242 ) );
  nand2 \comparator/C411  ( .a(\comparator/n807 ), .b(\comparator/n808 ), 
        .out(\comparator/N1240 ) );
  nand2 \comparator/C412  ( .a(\comparator/n809 ), .b(\comparator/n810 ), 
        .out(\comparator/N1238 ) );
  nand2 \comparator/C413  ( .a(\comparator/n811 ), .b(\comparator/n812 ), 
        .out(\comparator/N1236 ) );
  nand2 \comparator/C414  ( .a(\comparator/n813 ), .b(\comparator/n814 ), 
        .out(\comparator/N1234 ) );
  nand2 \comparator/C415  ( .a(\comparator/n815 ), .b(\comparator/n816 ), 
        .out(\comparator/N1232 ) );
  nand2 \comparator/C416  ( .a(\comparator/n817 ), .b(\comparator/n818 ), 
        .out(\comparator/N1230 ) );
  nand2 \comparator/C417  ( .a(\comparator/n819 ), .b(\comparator/n820 ), 
        .out(\comparator/N1228 ) );
  nand2 \comparator/C418  ( .a(\comparator/n821 ), .b(\comparator/n822 ), 
        .out(\comparator/N1226 ) );
  nand2 \comparator/C419  ( .a(\comparator/n823 ), .b(\comparator/n824 ), 
        .out(\comparator/N1224 ) );
  nand2 \comparator/C420  ( .a(\comparator/n825 ), .b(\comparator/n826 ), 
        .out(\comparator/N1222 ) );
  nand2 \comparator/C421  ( .a(\comparator/n827 ), .b(\comparator/n828 ), 
        .out(\comparator/N1220 ) );
  nand2 \comparator/C422  ( .a(\comparator/n829 ), .b(\comparator/n830 ), 
        .out(\comparator/N1218 ) );
  nand2 \comparator/C423  ( .a(\comparator/n831 ), .b(\comparator/n832 ), 
        .out(\comparator/N1216 ) );
  nand2 \comparator/C424  ( .a(\comparator/n833 ), .b(\comparator/n834 ), 
        .out(\comparator/N1214 ) );
  nand2 \comparator/C425  ( .a(\comparator/n835 ), .b(\comparator/n836 ), 
        .out(\comparator/N1212 ) );
  nand2 \comparator/C426  ( .a(\comparator/n837 ), .b(\comparator/n838 ), 
        .out(\comparator/N1210 ) );
  nand2 \comparator/C427  ( .a(\comparator/n839 ), .b(\comparator/n840 ), 
        .out(\comparator/N1208 ) );
  nand2 \comparator/C428  ( .a(\comparator/n841 ), .b(\comparator/n842 ), 
        .out(\comparator/N1206 ) );
  nand2 \comparator/C429  ( .a(\comparator/n843 ), .b(\comparator/n844 ), 
        .out(\comparator/N1204 ) );
  nand2 \comparator/C430  ( .a(\comparator/n845 ), .b(\comparator/n846 ), 
        .out(\comparator/N1202 ) );
  nand2 \comparator/C431  ( .a(\comparator/n847 ), .b(\comparator/n848 ), 
        .out(\comparator/N1200 ) );
  nand2 \comparator/C432  ( .a(\comparator/n849 ), .b(\comparator/n850 ), 
        .out(\comparator/N1198 ) );
  nand2 \comparator/C433  ( .a(\comparator/n851 ), .b(\comparator/n852 ), 
        .out(\comparator/N1196 ) );
  nand2 \comparator/C434  ( .a(\comparator/n853 ), .b(\comparator/n854 ), 
        .out(\comparator/N1194 ) );
  nand2 \comparator/C435  ( .a(\comparator/n855 ), .b(\comparator/n856 ), 
        .out(\comparator/N1192 ) );
  nand2 \comparator/C436  ( .a(\comparator/n857 ), .b(\comparator/n858 ), 
        .out(\comparator/N1190 ) );
  nand2 \comparator/C437  ( .a(\comparator/n859 ), .b(\comparator/n860 ), 
        .out(\comparator/N1188 ) );
  nand2 \comparator/C438  ( .a(\comparator/n861 ), .b(\comparator/n862 ), 
        .out(\comparator/N1186 ) );
  nand2 \comparator/C439  ( .a(\comparator/n863 ), .b(\comparator/n864 ), 
        .out(\comparator/N1184 ) );
  nand2 \comparator/C440  ( .a(\comparator/n865 ), .b(\comparator/n866 ), 
        .out(\comparator/N1182 ) );
  nand2 \comparator/C441  ( .a(\comparator/n867 ), .b(\comparator/n868 ), 
        .out(\comparator/N1180 ) );
  nand2 \comparator/C442  ( .a(\comparator/n869 ), .b(\comparator/n870 ), 
        .out(\comparator/N1178 ) );
  nand2 \comparator/C443  ( .a(\comparator/n871 ), .b(\comparator/n872 ), 
        .out(\comparator/N1176 ) );
  nand2 \comparator/C444  ( .a(\comparator/n873 ), .b(\comparator/n874 ), 
        .out(\comparator/N1174 ) );
  nand2 \comparator/C445  ( .a(\comparator/n875 ), .b(\comparator/n876 ), 
        .out(\comparator/N1172 ) );
  nand2 \comparator/C446  ( .a(\comparator/n877 ), .b(\comparator/n878 ), 
        .out(\comparator/N1170 ) );
  nand2 \comparator/C447  ( .a(\comparator/n879 ), .b(\comparator/n880 ), 
        .out(\comparator/N1168 ) );
  nand2 \comparator/C448  ( .a(\comparator/n881 ), .b(\comparator/n882 ), 
        .out(\comparator/N1166 ) );
  nand2 \comparator/C449  ( .a(\comparator/n883 ), .b(\comparator/n884 ), 
        .out(\comparator/N1164 ) );
  nand2 \comparator/C450  ( .a(\comparator/n885 ), .b(\comparator/n886 ), 
        .out(\comparator/N1162 ) );
  nand2 \comparator/C451  ( .a(\comparator/n887 ), .b(\comparator/n888 ), 
        .out(\comparator/N1160 ) );
  nand2 \comparator/C452  ( .a(\comparator/n889 ), .b(\comparator/n890 ), 
        .out(\comparator/N1158 ) );
  nand2 \comparator/C453  ( .a(\comparator/n891 ), .b(\comparator/n892 ), 
        .out(\comparator/N1156 ) );
  nand2 \comparator/C454  ( .a(\comparator/n893 ), .b(\comparator/n894 ), 
        .out(\comparator/N1154 ) );
  nand2 \comparator/C455  ( .a(\comparator/n895 ), .b(\comparator/n896 ), 
        .out(\comparator/N1152 ) );
  nand2 \comparator/C456  ( .a(\comparator/n897 ), .b(\comparator/n898 ), 
        .out(\comparator/N1150 ) );
  nand2 \comparator/C457  ( .a(\comparator/n899 ), .b(\comparator/n900 ), 
        .out(\comparator/N1148 ) );
  nand2 \comparator/C458  ( .a(\comparator/n901 ), .b(\comparator/n902 ), 
        .out(\comparator/N1146 ) );
  nand2 \comparator/C459  ( .a(\comparator/n903 ), .b(\comparator/n904 ), 
        .out(\comparator/N1144 ) );
  nand2 \comparator/C460  ( .a(\comparator/n905 ), .b(\comparator/n906 ), 
        .out(\comparator/N1142 ) );
  nand2 \comparator/C461  ( .a(\comparator/n907 ), .b(\comparator/n908 ), 
        .out(\comparator/N1140 ) );
  nand2 \comparator/C462  ( .a(\comparator/n909 ), .b(\comparator/n910 ), 
        .out(\comparator/N1138 ) );
  nand2 \comparator/C463  ( .a(\comparator/n911 ), .b(\comparator/n912 ), 
        .out(\comparator/N1136 ) );
  nand2 \comparator/C464  ( .a(\comparator/n913 ), .b(\comparator/n914 ), 
        .out(\comparator/N1134 ) );
  nand2 \comparator/C465  ( .a(\comparator/n915 ), .b(\comparator/n916 ), 
        .out(\comparator/N1132 ) );
  nand2 \comparator/C466  ( .a(\comparator/n917 ), .b(\comparator/n918 ), 
        .out(\comparator/N1130 ) );
  nand2 \comparator/C467  ( .a(\comparator/n919 ), .b(\comparator/n920 ), 
        .out(\comparator/N1128 ) );
  nand2 \comparator/C468  ( .a(\comparator/n921 ), .b(\comparator/n922 ), 
        .out(\comparator/N1126 ) );
  nand2 \comparator/C469  ( .a(\comparator/n923 ), .b(\comparator/n924 ), 
        .out(\comparator/N1124 ) );
  nand2 \comparator/C470  ( .a(\comparator/n925 ), .b(\comparator/n926 ), 
        .out(\comparator/N1122 ) );
  nand2 \comparator/C471  ( .a(\comparator/n927 ), .b(\comparator/n928 ), 
        .out(\comparator/N1120 ) );
  nand2 \comparator/C472  ( .a(\comparator/n929 ), .b(\comparator/n930 ), 
        .out(\comparator/N1118 ) );
  nand2 \comparator/C473  ( .a(\comparator/n931 ), .b(\comparator/n932 ), 
        .out(\comparator/N1116 ) );
  nand2 \comparator/C474  ( .a(\comparator/n933 ), .b(\comparator/n934 ), 
        .out(\comparator/N1114 ) );
  nand2 \comparator/C475  ( .a(\comparator/n935 ), .b(\comparator/n936 ), 
        .out(\comparator/N1112 ) );
  nand2 \comparator/C476  ( .a(\comparator/n937 ), .b(\comparator/n938 ), 
        .out(\comparator/N1110 ) );
  nand2 \comparator/C477  ( .a(\comparator/n939 ), .b(\comparator/n940 ), 
        .out(\comparator/N1108 ) );
  nand2 \comparator/C478  ( .a(\comparator/n941 ), .b(\comparator/n942 ), 
        .out(\comparator/N1106 ) );
  nand2 \comparator/C479  ( .a(\comparator/n943 ), .b(\comparator/n944 ), 
        .out(\comparator/N1104 ) );
  nand2 \comparator/C480  ( .a(\comparator/n945 ), .b(\comparator/n946 ), 
        .out(\comparator/N1102 ) );
  nand2 \comparator/C481  ( .a(\comparator/n947 ), .b(\comparator/n948 ), 
        .out(\comparator/N1100 ) );
  nand2 \comparator/C482  ( .a(\comparator/n949 ), .b(\comparator/n950 ), 
        .out(\comparator/N1098 ) );
  nand2 \comparator/C483  ( .a(\comparator/n951 ), .b(\comparator/n952 ), 
        .out(\comparator/N1096 ) );
  nand2 \comparator/C484  ( .a(\comparator/n953 ), .b(\comparator/n954 ), 
        .out(\comparator/N1094 ) );
  nand2 \comparator/C485  ( .a(\comparator/n955 ), .b(\comparator/n956 ), 
        .out(\comparator/N1092 ) );
  nand2 \comparator/C486  ( .a(\comparator/n957 ), .b(\comparator/n958 ), 
        .out(\comparator/N1090 ) );
  nand2 \comparator/C487  ( .a(\comparator/n959 ), .b(\comparator/n960 ), 
        .out(\comparator/N1088 ) );
  nand2 \comparator/C488  ( .a(\comparator/n961 ), .b(\comparator/n962 ), 
        .out(\comparator/N1086 ) );
  nand2 \comparator/C489  ( .a(\comparator/n963 ), .b(\comparator/n964 ), 
        .out(\comparator/N1084 ) );
  nand2 \comparator/C490  ( .a(\comparator/n965 ), .b(\comparator/n966 ), 
        .out(\comparator/N1082 ) );
  nand2 \comparator/C491  ( .a(\comparator/n967 ), .b(\comparator/n968 ), 
        .out(\comparator/N1080 ) );
  nand2 \comparator/C492  ( .a(\comparator/n969 ), .b(\comparator/n970 ), 
        .out(\comparator/N1078 ) );
  nand2 \comparator/C493  ( .a(\comparator/n971 ), .b(\comparator/n972 ), 
        .out(\comparator/N1076 ) );
  nand2 \comparator/C494  ( .a(\comparator/n973 ), .b(\comparator/n974 ), 
        .out(\comparator/N1074 ) );
  nand2 \comparator/C495  ( .a(\comparator/n975 ), .b(\comparator/n976 ), 
        .out(\comparator/N1072 ) );
  nand2 \comparator/C496  ( .a(\comparator/n977 ), .b(\comparator/n978 ), 
        .out(\comparator/N1070 ) );
  nand2 \comparator/C497  ( .a(\comparator/n979 ), .b(\comparator/n980 ), 
        .out(\comparator/N1068 ) );
  nand2 \comparator/C498  ( .a(\comparator/n981 ), .b(\comparator/n982 ), 
        .out(\comparator/N1066 ) );
  nand2 \comparator/C499  ( .a(\comparator/n983 ), .b(\comparator/n984 ), 
        .out(\comparator/N1064 ) );
  nand2 \comparator/C500  ( .a(\comparator/n985 ), .b(\comparator/n986 ), 
        .out(\comparator/N1062 ) );
  nand2 \comparator/C501  ( .a(\comparator/n987 ), .b(\comparator/n988 ), 
        .out(\comparator/N1060 ) );
  nand2 \comparator/C502  ( .a(\comparator/n989 ), .b(\comparator/n990 ), 
        .out(\comparator/N1058 ) );
  nand2 \comparator/C503  ( .a(\comparator/n991 ), .b(\comparator/n992 ), 
        .out(\comparator/N1056 ) );
  nand2 \comparator/C504  ( .a(\comparator/n993 ), .b(\comparator/n994 ), 
        .out(\comparator/N1054 ) );
  nand2 \comparator/C505  ( .a(\comparator/n995 ), .b(\comparator/n996 ), 
        .out(\comparator/N1052 ) );
  nand2 \comparator/C506  ( .a(\comparator/n997 ), .b(\comparator/n998 ), 
        .out(\comparator/N1050 ) );
  nand2 \comparator/C507  ( .a(\comparator/n999 ), .b(\comparator/n1000 ), 
        .out(\comparator/N1048 ) );
  nand2 \comparator/C508  ( .a(\comparator/n1001 ), .b(\comparator/n1002 ), 
        .out(\comparator/N1046 ) );
  nand2 \comparator/C509  ( .a(\comparator/n1003 ), .b(\comparator/n1004 ), 
        .out(\comparator/N1044 ) );
  nand2 \comparator/C510  ( .a(\comparator/n1005 ), .b(\comparator/n1006 ), 
        .out(\comparator/N1042 ) );
  nand2 \comparator/C511  ( .a(\comparator/n1007 ), .b(\comparator/n1008 ), 
        .out(\comparator/N1040 ) );
  nand2 \comparator/C512  ( .a(\comparator/n1009 ), .b(\comparator/n1010 ), 
        .out(\comparator/N1038 ) );
  nand2 \comparator/C513  ( .a(\comparator/n1011 ), .b(\comparator/n1012 ), 
        .out(\comparator/N1036 ) );
  nand2 \comparator/C514  ( .a(\comparator/n1013 ), .b(\comparator/n1014 ), 
        .out(\comparator/N1034 ) );
  nand2 \comparator/C515  ( .a(\comparator/n1015 ), .b(\comparator/n1016 ), 
        .out(\comparator/N1032 ) );
  nand2 \comparator/C516  ( .a(\comparator/n1017 ), .b(\comparator/n1018 ), 
        .out(\comparator/N1030 ) );
  nand2 \comparator/C517  ( .a(\comparator/n1019 ), .b(\comparator/n1020 ), 
        .out(\comparator/N1028 ) );
  nand2 \comparator/C518  ( .a(\comparator/n1021 ), .b(\comparator/n1022 ), 
        .out(\comparator/N1026 ) );
  nand2 \comparator/C519  ( .a(\comparator/n1023 ), .b(\comparator/n1024 ), 
        .out(\comparator/N1024 ) );
  nand2 \comparator/C520  ( .a(\comparator/n1025 ), .b(\comparator/n1026 ), 
        .out(\comparator/N1022 ) );
  nand2 \comparator/C521  ( .a(\comparator/n1027 ), .b(\comparator/n1028 ), 
        .out(\comparator/N1020 ) );
  nand2 \comparator/C522  ( .a(\comparator/n1029 ), .b(\comparator/n1030 ), 
        .out(\comparator/N1018 ) );
  nand2 \comparator/C523  ( .a(\comparator/n1031 ), .b(\comparator/n1032 ), 
        .out(\comparator/N1016 ) );
  nand2 \comparator/C524  ( .a(\comparator/n1033 ), .b(\comparator/n1034 ), 
        .out(\comparator/N1014 ) );
  nand2 \comparator/C525  ( .a(\comparator/n1035 ), .b(\comparator/n1036 ), 
        .out(\comparator/N1012 ) );
  nand2 \comparator/C526  ( .a(\comparator/n1037 ), .b(\comparator/n1038 ), 
        .out(\comparator/N1010 ) );
  nand2 \comparator/C527  ( .a(\comparator/n1039 ), .b(\comparator/n1040 ), 
        .out(\comparator/N1008 ) );
  nand2 \comparator/C528  ( .a(\comparator/n1041 ), .b(\comparator/n1042 ), 
        .out(\comparator/N1006 ) );
  nand2 \comparator/C529  ( .a(\comparator/n1043 ), .b(\comparator/n1044 ), 
        .out(\comparator/N1004 ) );
  nand2 \comparator/C530  ( .a(\comparator/n1045 ), .b(\comparator/n1046 ), 
        .out(\comparator/N1002 ) );
  nand2 \comparator/C531  ( .a(\comparator/n1047 ), .b(\comparator/n1048 ), 
        .out(\comparator/N1000 ) );
  nand2 \comparator/C532  ( .a(\comparator/n1049 ), .b(\comparator/n1050 ), 
        .out(\comparator/N998 ) );
  nand2 \comparator/C533  ( .a(\comparator/n1051 ), .b(\comparator/n1052 ), 
        .out(\comparator/N996 ) );
  nand2 \comparator/C534  ( .a(\comparator/n1053 ), .b(\comparator/n1054 ), 
        .out(\comparator/N994 ) );
  nand2 \comparator/C535  ( .a(\comparator/n1055 ), .b(\comparator/n1056 ), 
        .out(\comparator/N992 ) );
  nand2 \comparator/C536  ( .a(\comparator/n1057 ), .b(\comparator/n1058 ), 
        .out(\comparator/N990 ) );
  nand2 \comparator/C537  ( .a(\comparator/n1059 ), .b(\comparator/n1060 ), 
        .out(\comparator/N988 ) );
  nand2 \comparator/C538  ( .a(\comparator/n1061 ), .b(\comparator/n1062 ), 
        .out(\comparator/N986 ) );
  nand2 \comparator/C539  ( .a(\comparator/n1063 ), .b(\comparator/n1064 ), 
        .out(\comparator/N984 ) );
  nand2 \comparator/C540  ( .a(\comparator/n1065 ), .b(\comparator/n1066 ), 
        .out(\comparator/N982 ) );
  nand2 \comparator/C541  ( .a(\comparator/n1067 ), .b(\comparator/n1068 ), 
        .out(\comparator/N980 ) );
  nand2 \comparator/C542  ( .a(\comparator/n1069 ), .b(\comparator/n1070 ), 
        .out(\comparator/N978 ) );
  nand2 \comparator/C543  ( .a(\comparator/n1071 ), .b(\comparator/n1072 ), 
        .out(\comparator/N976 ) );
  nand2 \comparator/C544  ( .a(\comparator/n1073 ), .b(\comparator/n1074 ), 
        .out(\comparator/N974 ) );
  nand2 \comparator/C545  ( .a(\comparator/n1075 ), .b(\comparator/n1076 ), 
        .out(\comparator/N972 ) );
  nand2 \comparator/C546  ( .a(\comparator/n1077 ), .b(\comparator/n1078 ), 
        .out(\comparator/N970 ) );
  nand2 \comparator/C547  ( .a(\comparator/n1079 ), .b(\comparator/n1080 ), 
        .out(\comparator/N968 ) );
  nand2 \comparator/C548  ( .a(\comparator/n1081 ), .b(\comparator/n1082 ), 
        .out(\comparator/N966 ) );
  nand2 \comparator/C549  ( .a(\comparator/n1083 ), .b(\comparator/n1084 ), 
        .out(\comparator/N964 ) );
  nand2 \comparator/C550  ( .a(\comparator/n1085 ), .b(\comparator/n1086 ), 
        .out(\comparator/N962 ) );
  nand2 \comparator/C551  ( .a(\comparator/n1087 ), .b(\comparator/n1088 ), 
        .out(\comparator/N960 ) );
  nand2 \comparator/C552  ( .a(\comparator/n1089 ), .b(\comparator/n1090 ), 
        .out(\comparator/N958 ) );
  nand2 \comparator/C553  ( .a(\comparator/n1091 ), .b(\comparator/n1092 ), 
        .out(\comparator/N956 ) );
  nand2 \comparator/C554  ( .a(\comparator/n1093 ), .b(\comparator/n1094 ), 
        .out(\comparator/N954 ) );
  nand2 \comparator/C555  ( .a(\comparator/n1095 ), .b(\comparator/n1096 ), 
        .out(\comparator/N952 ) );
  nand2 \comparator/C556  ( .a(\comparator/n1097 ), .b(\comparator/n1098 ), 
        .out(\comparator/N950 ) );
  nand2 \comparator/C557  ( .a(\comparator/n1099 ), .b(\comparator/n1100 ), 
        .out(\comparator/N948 ) );
  nand2 \comparator/C558  ( .a(\comparator/n1101 ), .b(\comparator/n1102 ), 
        .out(\comparator/N946 ) );
  nand2 \comparator/C559  ( .a(\comparator/n1103 ), .b(\comparator/n1104 ), 
        .out(\comparator/N944 ) );
  nand2 \comparator/C560  ( .a(\comparator/n1105 ), .b(\comparator/n1106 ), 
        .out(\comparator/N942 ) );
  nand2 \comparator/C561  ( .a(\comparator/n1107 ), .b(\comparator/n1108 ), 
        .out(\comparator/N940 ) );
  nand2 \comparator/C562  ( .a(\comparator/n1109 ), .b(\comparator/n1110 ), 
        .out(\comparator/N938 ) );
  nand2 \comparator/C563  ( .a(\comparator/n1111 ), .b(\comparator/n1112 ), 
        .out(\comparator/N936 ) );
  nand2 \comparator/C564  ( .a(\comparator/n1113 ), .b(\comparator/n1114 ), 
        .out(\comparator/N934 ) );
  nand2 \comparator/C565  ( .a(\comparator/n1115 ), .b(\comparator/n1116 ), 
        .out(\comparator/N932 ) );
  nand2 \comparator/C566  ( .a(\comparator/n1117 ), .b(\comparator/n1118 ), 
        .out(\comparator/N930 ) );
  nand2 \comparator/C567  ( .a(\comparator/n1119 ), .b(\comparator/n1120 ), 
        .out(\comparator/N928 ) );
  nand2 \comparator/C568  ( .a(\comparator/n1121 ), .b(\comparator/n1122 ), 
        .out(\comparator/N926 ) );
  nand2 \comparator/C569  ( .a(\comparator/n1123 ), .b(\comparator/n1124 ), 
        .out(\comparator/N924 ) );
  nand2 \comparator/C570  ( .a(\comparator/n1125 ), .b(\comparator/n1126 ), 
        .out(\comparator/N922 ) );
  nand2 \comparator/C571  ( .a(\comparator/n1127 ), .b(\comparator/n1128 ), 
        .out(\comparator/N920 ) );
  nand2 \comparator/C572  ( .a(\comparator/n1129 ), .b(\comparator/n1130 ), 
        .out(\comparator/N918 ) );
  nand2 \comparator/C573  ( .a(\comparator/n1131 ), .b(\comparator/n1132 ), 
        .out(\comparator/N916 ) );
  nand2 \comparator/C574  ( .a(\comparator/n1133 ), .b(\comparator/n1134 ), 
        .out(\comparator/N914 ) );
  nand2 \comparator/C575  ( .a(\comparator/n1135 ), .b(\comparator/n1136 ), 
        .out(\comparator/N912 ) );
  nand2 \comparator/C576  ( .a(\comparator/n1137 ), .b(\comparator/n1138 ), 
        .out(\comparator/N910 ) );
  nand2 \comparator/C577  ( .a(\comparator/n1139 ), .b(\comparator/n1140 ), 
        .out(\comparator/N908 ) );
  nand2 \comparator/C578  ( .a(\comparator/n1141 ), .b(\comparator/n1142 ), 
        .out(\comparator/N906 ) );
  nand2 \comparator/C579  ( .a(\comparator/n1143 ), .b(\comparator/n1144 ), 
        .out(\comparator/N904 ) );
  nand2 \comparator/C580  ( .a(\comparator/n1145 ), .b(\comparator/n1146 ), 
        .out(\comparator/N902 ) );
  nand2 \comparator/C581  ( .a(\comparator/n1147 ), .b(\comparator/n1148 ), 
        .out(\comparator/N900 ) );
  nand2 \comparator/C582  ( .a(\comparator/n1149 ), .b(\comparator/n1150 ), 
        .out(\comparator/N898 ) );
  nand2 \comparator/C583  ( .a(\comparator/n1151 ), .b(\comparator/n1152 ), 
        .out(\comparator/N896 ) );
  nand2 \comparator/C584  ( .a(\comparator/n1153 ), .b(\comparator/n1154 ), 
        .out(\comparator/N894 ) );
  nand2 \comparator/C585  ( .a(\comparator/n1155 ), .b(\comparator/n1156 ), 
        .out(\comparator/N892 ) );
  nand2 \comparator/C586  ( .a(\comparator/n1157 ), .b(\comparator/n1158 ), 
        .out(\comparator/N890 ) );
  nand2 \comparator/C587  ( .a(\comparator/n1159 ), .b(\comparator/n1160 ), 
        .out(\comparator/N888 ) );
  nand2 \comparator/C588  ( .a(\comparator/n1161 ), .b(\comparator/n1162 ), 
        .out(\comparator/N886 ) );
  nand2 \comparator/C589  ( .a(\comparator/n1163 ), .b(\comparator/n1164 ), 
        .out(\comparator/N884 ) );
  nand2 \comparator/C590  ( .a(\comparator/n1165 ), .b(\comparator/n1166 ), 
        .out(\comparator/N882 ) );
  nand2 \comparator/C591  ( .a(\comparator/n1167 ), .b(\comparator/n1168 ), 
        .out(\comparator/N880 ) );
  nand2 \comparator/C592  ( .a(\comparator/n1169 ), .b(\comparator/n1170 ), 
        .out(\comparator/N878 ) );
  nand2 \comparator/C593  ( .a(\comparator/n1171 ), .b(\comparator/n1172 ), 
        .out(\comparator/N876 ) );
  nand2 \comparator/C594  ( .a(\comparator/n1173 ), .b(\comparator/n1174 ), 
        .out(\comparator/N874 ) );
  nand2 \comparator/C595  ( .a(\comparator/n1175 ), .b(\comparator/n1176 ), 
        .out(\comparator/N872 ) );
  nand2 \comparator/C596  ( .a(\comparator/n1177 ), .b(\comparator/n1178 ), 
        .out(\comparator/N870 ) );
  nand2 \comparator/C597  ( .a(\comparator/n1179 ), .b(\comparator/n1180 ), 
        .out(\comparator/N868 ) );
  nand2 \comparator/C598  ( .a(\comparator/n1181 ), .b(\comparator/n1182 ), 
        .out(\comparator/N866 ) );
  nand2 \comparator/C599  ( .a(\comparator/n1183 ), .b(\comparator/n1184 ), 
        .out(\comparator/N864 ) );
  nand2 \comparator/C600  ( .a(\comparator/n1185 ), .b(\comparator/n1186 ), 
        .out(\comparator/N862 ) );
  nand2 \comparator/C601  ( .a(\comparator/n1187 ), .b(\comparator/n1188 ), 
        .out(\comparator/N860 ) );
  nand2 \comparator/C602  ( .a(\comparator/n1189 ), .b(\comparator/n1190 ), 
        .out(\comparator/N858 ) );
  nand2 \comparator/C603  ( .a(\comparator/n1191 ), .b(\comparator/n1192 ), 
        .out(\comparator/N856 ) );
  nand2 \comparator/C604  ( .a(\comparator/n1193 ), .b(\comparator/n1194 ), 
        .out(\comparator/N854 ) );
  nand2 \comparator/C605  ( .a(\comparator/n1195 ), .b(\comparator/n1196 ), 
        .out(\comparator/N852 ) );
  nand2 \comparator/C606  ( .a(\comparator/n1197 ), .b(\comparator/n1198 ), 
        .out(\comparator/N850 ) );
  nand2 \comparator/C607  ( .a(\comparator/n1199 ), .b(\comparator/n1200 ), 
        .out(\comparator/N848 ) );
  nand2 \comparator/C608  ( .a(\comparator/n1201 ), .b(\comparator/n1202 ), 
        .out(\comparator/N846 ) );
  nand2 \comparator/C609  ( .a(\comparator/n1203 ), .b(\comparator/n1204 ), 
        .out(\comparator/N844 ) );
  nand2 \comparator/C610  ( .a(\comparator/n1205 ), .b(\comparator/n1206 ), 
        .out(\comparator/N842 ) );
  nand2 \comparator/C611  ( .a(\comparator/n1207 ), .b(\comparator/n1208 ), 
        .out(\comparator/N840 ) );
  nand2 \comparator/C612  ( .a(\comparator/n1209 ), .b(\comparator/n1210 ), 
        .out(\comparator/N838 ) );
  nand2 \comparator/C613  ( .a(\comparator/n1211 ), .b(\comparator/n1212 ), 
        .out(\comparator/N836 ) );
  nand2 \comparator/C614  ( .a(\comparator/n1213 ), .b(\comparator/n1214 ), 
        .out(\comparator/N834 ) );
  nand2 \comparator/C615  ( .a(\comparator/n1215 ), .b(\comparator/n1216 ), 
        .out(\comparator/N832 ) );
  nand2 \comparator/C616  ( .a(\comparator/n1217 ), .b(\comparator/n1218 ), 
        .out(\comparator/N830 ) );
  nand2 \comparator/C617  ( .a(\comparator/n1219 ), .b(\comparator/n1220 ), 
        .out(\comparator/N828 ) );
  nand2 \comparator/C618  ( .a(\comparator/n1221 ), .b(\comparator/n1222 ), 
        .out(\comparator/N826 ) );
  nand2 \comparator/C619  ( .a(\comparator/n1223 ), .b(\comparator/n1224 ), 
        .out(\comparator/N824 ) );
  nand2 \comparator/C620  ( .a(\comparator/n1225 ), .b(\comparator/n1226 ), 
        .out(\comparator/N822 ) );
  nand2 \comparator/C621  ( .a(\comparator/n1227 ), .b(\comparator/n1228 ), 
        .out(\comparator/N820 ) );
  nand2 \comparator/C622  ( .a(\comparator/n1229 ), .b(\comparator/n1230 ), 
        .out(\comparator/N818 ) );
  nand2 \comparator/C623  ( .a(\comparator/n1231 ), .b(\comparator/n1232 ), 
        .out(\comparator/N816 ) );
  nand2 \comparator/C624  ( .a(\comparator/n1233 ), .b(\comparator/n1234 ), 
        .out(\comparator/N814 ) );
  nand2 \comparator/C625  ( .a(\comparator/n1235 ), .b(\comparator/n1236 ), 
        .out(\comparator/N812 ) );
  nand2 \comparator/C626  ( .a(\comparator/n1237 ), .b(\comparator/n1238 ), 
        .out(\comparator/N810 ) );
  nand2 \comparator/C627  ( .a(\comparator/n1239 ), .b(\comparator/n1240 ), 
        .out(\comparator/N808 ) );
  nand2 \comparator/C628  ( .a(\comparator/n1241 ), .b(\comparator/n1242 ), 
        .out(\comparator/N806 ) );
  nand2 \comparator/C629  ( .a(\comparator/n1243 ), .b(\comparator/n1244 ), 
        .out(\comparator/N804 ) );
  nand2 \comparator/C630  ( .a(\comparator/n1245 ), .b(\comparator/n1246 ), 
        .out(\comparator/N802 ) );
  nand2 \comparator/C631  ( .a(\comparator/n1247 ), .b(\comparator/n1248 ), 
        .out(\comparator/N800 ) );
  nand2 \comparator/C632  ( .a(\comparator/n1249 ), .b(\comparator/n1250 ), 
        .out(\comparator/N798 ) );
  nand2 \comparator/C633  ( .a(\comparator/n1251 ), .b(\comparator/n1252 ), 
        .out(\comparator/N796 ) );
  nand2 \comparator/C634  ( .a(\comparator/n1253 ), .b(\comparator/n1254 ), 
        .out(\comparator/N794 ) );
  nand2 \comparator/C635  ( .a(\comparator/n1255 ), .b(\comparator/n1256 ), 
        .out(\comparator/N792 ) );
  nand2 \comparator/C636  ( .a(\comparator/n1257 ), .b(\comparator/n1258 ), 
        .out(\comparator/N790 ) );
  nand2 \comparator/C637  ( .a(\comparator/n1259 ), .b(\comparator/n1260 ), 
        .out(\comparator/N788 ) );
  nand2 \comparator/C638  ( .a(\comparator/n1261 ), .b(\comparator/n1262 ), 
        .out(\comparator/N786 ) );
  nand2 \comparator/C639  ( .a(\comparator/n1263 ), .b(\comparator/n1264 ), 
        .out(\comparator/N784 ) );
  nand2 \comparator/C640  ( .a(\comparator/n1265 ), .b(\comparator/n1266 ), 
        .out(\comparator/N782 ) );
  nand2 \comparator/C641  ( .a(\comparator/n1267 ), .b(\comparator/n1268 ), 
        .out(\comparator/N780 ) );
  nand2 \comparator/C642  ( .a(\comparator/n1269 ), .b(\comparator/n1270 ), 
        .out(\comparator/N778 ) );
  nand2 \comparator/C643  ( .a(\comparator/n1271 ), .b(\comparator/n1272 ), 
        .out(\comparator/N776 ) );
  nand2 \comparator/C644  ( .a(\comparator/n1273 ), .b(\comparator/n1274 ), 
        .out(\comparator/N774 ) );
  nand2 \comparator/C645  ( .a(\comparator/n1275 ), .b(\comparator/n1276 ), 
        .out(\comparator/N772 ) );
  nand2 \comparator/C646  ( .a(\comparator/n1277 ), .b(\comparator/n1278 ), 
        .out(\comparator/N770 ) );
  nand2 \comparator/C647  ( .a(\comparator/n1279 ), .b(\comparator/n1280 ), 
        .out(\comparator/N768 ) );
  nand2 \comparator/C648  ( .a(\comparator/n1281 ), .b(\comparator/n1282 ), 
        .out(\comparator/N766 ) );
  nand2 \comparator/C649  ( .a(\comparator/n1283 ), .b(\comparator/n1284 ), 
        .out(\comparator/N764 ) );
  nand2 \comparator/C650  ( .a(\comparator/n1285 ), .b(\comparator/n1286 ), 
        .out(\comparator/N762 ) );
  nand2 \comparator/C651  ( .a(\comparator/n1287 ), .b(\comparator/n1288 ), 
        .out(\comparator/N760 ) );
  nand2 \comparator/C652  ( .a(\comparator/n1289 ), .b(\comparator/n1290 ), 
        .out(\comparator/N758 ) );
  nand2 \comparator/C653  ( .a(\comparator/n1291 ), .b(\comparator/n1292 ), 
        .out(\comparator/N756 ) );
  nand2 \comparator/C654  ( .a(\comparator/n1293 ), .b(\comparator/n1294 ), 
        .out(\comparator/N754 ) );
  nand2 \comparator/C655  ( .a(\comparator/n1295 ), .b(\comparator/n1296 ), 
        .out(\comparator/N752 ) );
  nand2 \comparator/C656  ( .a(\comparator/n1297 ), .b(\comparator/n1298 ), 
        .out(\comparator/N750 ) );
  nand2 \comparator/C657  ( .a(\comparator/n1299 ), .b(\comparator/n1300 ), 
        .out(\comparator/N748 ) );
  nand2 \comparator/C658  ( .a(\comparator/n1301 ), .b(\comparator/n1302 ), 
        .out(\comparator/N746 ) );
  nand2 \comparator/C659  ( .a(\comparator/n1303 ), .b(\comparator/n1304 ), 
        .out(\comparator/N744 ) );
  nand2 \comparator/C660  ( .a(\comparator/n1305 ), .b(\comparator/n1306 ), 
        .out(\comparator/N742 ) );
  nand2 \comparator/C661  ( .a(\comparator/n1307 ), .b(\comparator/n1308 ), 
        .out(\comparator/N740 ) );
  nand2 \comparator/C662  ( .a(\comparator/n1309 ), .b(\comparator/n1310 ), 
        .out(\comparator/N738 ) );
  nand2 \comparator/C663  ( .a(\comparator/n1311 ), .b(\comparator/n1312 ), 
        .out(\comparator/N736 ) );
  nand2 \comparator/C664  ( .a(\comparator/n1313 ), .b(\comparator/n1314 ), 
        .out(\comparator/N734 ) );
  nand2 \comparator/C665  ( .a(\comparator/n1315 ), .b(\comparator/n1316 ), 
        .out(\comparator/N732 ) );
  nand2 \comparator/C666  ( .a(\comparator/n1317 ), .b(\comparator/n1318 ), 
        .out(\comparator/N730 ) );
  nand2 \comparator/C667  ( .a(\comparator/n1319 ), .b(\comparator/n1320 ), 
        .out(\comparator/N728 ) );
  nand2 \comparator/C668  ( .a(\comparator/n1321 ), .b(\comparator/n1322 ), 
        .out(\comparator/N726 ) );
  nand2 \comparator/C669  ( .a(\comparator/n1323 ), .b(\comparator/n1324 ), 
        .out(\comparator/N724 ) );
  nand2 \comparator/C670  ( .a(\comparator/n1325 ), .b(\comparator/n1326 ), 
        .out(\comparator/N722 ) );
  nand2 \comparator/C671  ( .a(\comparator/n1327 ), .b(\comparator/n1328 ), 
        .out(\comparator/N720 ) );
  nand2 \comparator/C672  ( .a(\comparator/n1329 ), .b(\comparator/n1330 ), 
        .out(\comparator/N718 ) );
  nand2 \comparator/C673  ( .a(\comparator/n1331 ), .b(\comparator/n1332 ), 
        .out(\comparator/N716 ) );
  nand2 \comparator/C674  ( .a(\comparator/n1333 ), .b(\comparator/n1334 ), 
        .out(\comparator/N714 ) );
  nand2 \comparator/C675  ( .a(\comparator/n1335 ), .b(\comparator/n1336 ), 
        .out(\comparator/N712 ) );
  nand2 \comparator/C676  ( .a(\comparator/n1337 ), .b(\comparator/n1338 ), 
        .out(\comparator/N710 ) );
  nand2 \comparator/C677  ( .a(\comparator/n1339 ), .b(\comparator/n1340 ), 
        .out(\comparator/N708 ) );
  nand2 \comparator/C678  ( .a(\comparator/n1341 ), .b(\comparator/n1342 ), 
        .out(\comparator/N706 ) );
  nand2 \comparator/C679  ( .a(\comparator/n1343 ), .b(\comparator/n1344 ), 
        .out(\comparator/N704 ) );
  nand2 \comparator/C680  ( .a(\comparator/n1345 ), .b(\comparator/n1346 ), 
        .out(\comparator/N702 ) );
  nand2 \comparator/C681  ( .a(\comparator/n1347 ), .b(\comparator/n1348 ), 
        .out(\comparator/N700 ) );
  nand2 \comparator/C682  ( .a(\comparator/n1349 ), .b(\comparator/n1350 ), 
        .out(\comparator/N698 ) );
  nand2 \comparator/C683  ( .a(\comparator/n1351 ), .b(\comparator/n1352 ), 
        .out(\comparator/N696 ) );
  nand2 \comparator/C684  ( .a(\comparator/n1353 ), .b(\comparator/n1354 ), 
        .out(\comparator/N694 ) );
  nand2 \comparator/C685  ( .a(\comparator/n1355 ), .b(\comparator/n1356 ), 
        .out(\comparator/N692 ) );
  nand2 \comparator/C686  ( .a(\comparator/n1357 ), .b(\comparator/n1358 ), 
        .out(\comparator/N690 ) );
  nand2 \comparator/C687  ( .a(\comparator/n1359 ), .b(\comparator/n1360 ), 
        .out(\comparator/N688 ) );
  nand2 \comparator/C688  ( .a(\comparator/n1361 ), .b(\comparator/n1362 ), 
        .out(\comparator/N686 ) );
  nand2 \comparator/C689  ( .a(\comparator/n1363 ), .b(\comparator/n1364 ), 
        .out(\comparator/N684 ) );
  nand2 \comparator/C690  ( .a(\comparator/n1365 ), .b(\comparator/n1366 ), 
        .out(\comparator/N682 ) );
  nand2 \comparator/C691  ( .a(\comparator/n1367 ), .b(\comparator/n1368 ), 
        .out(\comparator/N680 ) );
  nand2 \comparator/C692  ( .a(\comparator/n1369 ), .b(\comparator/n1370 ), 
        .out(\comparator/N678 ) );
  nand2 \comparator/C693  ( .a(\comparator/n1371 ), .b(\comparator/n1372 ), 
        .out(\comparator/N676 ) );
  nand2 \comparator/C694  ( .a(\comparator/n1373 ), .b(\comparator/n1374 ), 
        .out(\comparator/N674 ) );
  nand2 \comparator/C695  ( .a(\comparator/n1375 ), .b(\comparator/n1376 ), 
        .out(\comparator/N672 ) );
  nand2 \comparator/C696  ( .a(\comparator/n1377 ), .b(\comparator/n1378 ), 
        .out(\comparator/N670 ) );
  nand2 \comparator/C697  ( .a(\comparator/n1379 ), .b(\comparator/n1380 ), 
        .out(\comparator/N668 ) );
  nand2 \comparator/C698  ( .a(\comparator/n1381 ), .b(\comparator/n1382 ), 
        .out(\comparator/N666 ) );
  nand2 \comparator/C699  ( .a(\comparator/n1383 ), .b(\comparator/n1384 ), 
        .out(\comparator/N664 ) );
  nand2 \comparator/C700  ( .a(\comparator/n1385 ), .b(\comparator/n1386 ), 
        .out(\comparator/N662 ) );
  nand2 \comparator/C701  ( .a(\comparator/n1387 ), .b(\comparator/n1388 ), 
        .out(\comparator/N660 ) );
  nand2 \comparator/C702  ( .a(\comparator/n1389 ), .b(\comparator/n1390 ), 
        .out(\comparator/N658 ) );
  nand2 \comparator/C703  ( .a(\comparator/n1391 ), .b(\comparator/n1392 ), 
        .out(\comparator/N656 ) );
  nand2 \comparator/C704  ( .a(\comparator/n1393 ), .b(\comparator/n1394 ), 
        .out(\comparator/N654 ) );
  nand2 \comparator/C705  ( .a(\comparator/n1395 ), .b(\comparator/n1396 ), 
        .out(\comparator/N652 ) );
  nand2 \comparator/C706  ( .a(\comparator/n1397 ), .b(\comparator/n1398 ), 
        .out(\comparator/N650 ) );
  nand2 \comparator/C707  ( .a(\comparator/n1399 ), .b(\comparator/n1400 ), 
        .out(\comparator/N648 ) );
  nand2 \comparator/C708  ( .a(\comparator/n1401 ), .b(\comparator/n1402 ), 
        .out(\comparator/N646 ) );
  nand2 \comparator/C709  ( .a(\comparator/n1403 ), .b(\comparator/n1404 ), 
        .out(\comparator/N644 ) );
  nand2 \comparator/C710  ( .a(\comparator/n1405 ), .b(\comparator/n1406 ), 
        .out(\comparator/N642 ) );
  nand2 \comparator/C711  ( .a(\comparator/n1407 ), .b(\comparator/n1408 ), 
        .out(\comparator/N640 ) );
  nand2 \comparator/C712  ( .a(\comparator/n1409 ), .b(\comparator/n1410 ), 
        .out(\comparator/N638 ) );
  nand2 \comparator/C713  ( .a(\comparator/n1411 ), .b(\comparator/n1412 ), 
        .out(\comparator/N636 ) );
  nand2 \comparator/C714  ( .a(\comparator/n1413 ), .b(\comparator/n1414 ), 
        .out(\comparator/N634 ) );
  nand2 \comparator/C715  ( .a(\comparator/n1415 ), .b(\comparator/n1416 ), 
        .out(\comparator/N632 ) );
  nand2 \comparator/C716  ( .a(\comparator/n1417 ), .b(\comparator/n1418 ), 
        .out(\comparator/N630 ) );
  nand2 \comparator/C717  ( .a(\comparator/n1419 ), .b(\comparator/n1420 ), 
        .out(\comparator/N628 ) );
  nand2 \comparator/C718  ( .a(\comparator/n1421 ), .b(\comparator/n1422 ), 
        .out(\comparator/N626 ) );
  nand2 \comparator/C719  ( .a(\comparator/n1423 ), .b(\comparator/n1424 ), 
        .out(\comparator/N624 ) );
  nand2 \comparator/C720  ( .a(\comparator/n1425 ), .b(\comparator/n1426 ), 
        .out(\comparator/N622 ) );
  nand2 \comparator/C721  ( .a(\comparator/n1427 ), .b(\comparator/n1428 ), 
        .out(\comparator/N620 ) );
  nand2 \comparator/C722  ( .a(\comparator/n1429 ), .b(\comparator/n1430 ), 
        .out(\comparator/N618 ) );
  nand2 \comparator/C723  ( .a(\comparator/n1431 ), .b(\comparator/n1432 ), 
        .out(\comparator/N616 ) );
  nand2 \comparator/C724  ( .a(\comparator/n1433 ), .b(\comparator/n1434 ), 
        .out(\comparator/N614 ) );
  nand2 \comparator/C725  ( .a(\comparator/n1435 ), .b(\comparator/n1436 ), 
        .out(\comparator/N612 ) );
  nand2 \comparator/C726  ( .a(\comparator/n1437 ), .b(\comparator/n1438 ), 
        .out(\comparator/N610 ) );
  nand2 \comparator/C727  ( .a(\comparator/n1439 ), .b(\comparator/n1440 ), 
        .out(\comparator/N608 ) );
  nand2 \comparator/C728  ( .a(\comparator/n1441 ), .b(\comparator/n1442 ), 
        .out(\comparator/N606 ) );
  nand2 \comparator/C729  ( .a(\comparator/n1443 ), .b(\comparator/n1444 ), 
        .out(\comparator/N604 ) );
  nand2 \comparator/C730  ( .a(\comparator/n1445 ), .b(\comparator/n1446 ), 
        .out(\comparator/N602 ) );
  nand2 \comparator/C731  ( .a(\comparator/n1447 ), .b(\comparator/n1448 ), 
        .out(\comparator/N600 ) );
  nand2 \comparator/C732  ( .a(\comparator/n1449 ), .b(\comparator/n1450 ), 
        .out(\comparator/N598 ) );
  nand2 \comparator/C733  ( .a(\comparator/n1451 ), .b(\comparator/n1452 ), 
        .out(\comparator/N596 ) );
  nand2 \comparator/C734  ( .a(\comparator/n1453 ), .b(\comparator/n1454 ), 
        .out(\comparator/N594 ) );
  nand2 \comparator/C735  ( .a(\comparator/n1455 ), .b(\comparator/n1456 ), 
        .out(\comparator/N592 ) );
  nand2 \comparator/C736  ( .a(\comparator/n1457 ), .b(\comparator/n1458 ), 
        .out(\comparator/N590 ) );
  nand2 \comparator/C737  ( .a(\comparator/n1459 ), .b(\comparator/n1460 ), 
        .out(\comparator/N588 ) );
  nand2 \comparator/C738  ( .a(\comparator/n1461 ), .b(\comparator/n1462 ), 
        .out(\comparator/N586 ) );
  nand2 \comparator/C739  ( .a(\comparator/n1463 ), .b(\comparator/n1464 ), 
        .out(\comparator/N584 ) );
  nand2 \comparator/C740  ( .a(\comparator/n1465 ), .b(\comparator/n1466 ), 
        .out(\comparator/N582 ) );
  nand2 \comparator/C741  ( .a(\comparator/n1467 ), .b(\comparator/n1468 ), 
        .out(\comparator/N580 ) );
  nand2 \comparator/C742  ( .a(\comparator/n1469 ), .b(\comparator/n1470 ), 
        .out(\comparator/N578 ) );
  nand2 \comparator/C743  ( .a(\comparator/n1471 ), .b(\comparator/n1472 ), 
        .out(\comparator/N576 ) );
  nand2 \comparator/C744  ( .a(\comparator/n1473 ), .b(\comparator/n1474 ), 
        .out(\comparator/N574 ) );
  nand2 \comparator/C745  ( .a(\comparator/n1475 ), .b(\comparator/n1476 ), 
        .out(\comparator/N572 ) );
  nand2 \comparator/C746  ( .a(\comparator/n1477 ), .b(\comparator/n1478 ), 
        .out(\comparator/N570 ) );
  nand2 \comparator/C747  ( .a(\comparator/n1479 ), .b(\comparator/n1480 ), 
        .out(\comparator/N568 ) );
  nand2 \comparator/C748  ( .a(\comparator/n1481 ), .b(\comparator/n1482 ), 
        .out(\comparator/N566 ) );
  nand2 \comparator/C749  ( .a(\comparator/n1483 ), .b(\comparator/n1484 ), 
        .out(\comparator/N564 ) );
  nand2 \comparator/C750  ( .a(\comparator/n1485 ), .b(\comparator/n1486 ), 
        .out(\comparator/N562 ) );
  nand2 \comparator/C751  ( .a(\comparator/n1487 ), .b(\comparator/n1488 ), 
        .out(\comparator/N560 ) );
  nand2 \comparator/C752  ( .a(\comparator/n1489 ), .b(\comparator/n1490 ), 
        .out(\comparator/N558 ) );
  nand2 \comparator/C753  ( .a(\comparator/n1491 ), .b(\comparator/n1492 ), 
        .out(\comparator/N556 ) );
  nand2 \comparator/C754  ( .a(\comparator/n1493 ), .b(\comparator/n1494 ), 
        .out(\comparator/N554 ) );
  nand2 \comparator/C755  ( .a(\comparator/n1495 ), .b(\comparator/n1496 ), 
        .out(\comparator/N552 ) );
  nand2 \comparator/C756  ( .a(\comparator/n1497 ), .b(\comparator/n1498 ), 
        .out(\comparator/N550 ) );
  nand2 \comparator/C757  ( .a(\comparator/n1499 ), .b(\comparator/n1500 ), 
        .out(\comparator/N548 ) );
  nand2 \comparator/C758  ( .a(\comparator/n1501 ), .b(\comparator/n1502 ), 
        .out(\comparator/N546 ) );
  nand2 \comparator/C759  ( .a(\comparator/n1503 ), .b(\comparator/n1504 ), 
        .out(\comparator/N544 ) );
  nand2 \comparator/C760  ( .a(\comparator/n1505 ), .b(\comparator/n1506 ), 
        .out(\comparator/N542 ) );
  nand2 \comparator/C761  ( .a(\comparator/n1507 ), .b(\comparator/n1508 ), 
        .out(\comparator/N540 ) );
  nand2 \comparator/C762  ( .a(\comparator/n1509 ), .b(\comparator/n1510 ), 
        .out(\comparator/N538 ) );
  nand2 \comparator/C763  ( .a(\comparator/n1511 ), .b(\comparator/n1512 ), 
        .out(\comparator/N536 ) );
  nand2 \comparator/C764  ( .a(\comparator/n1513 ), .b(\comparator/n1514 ), 
        .out(\comparator/N534 ) );
  nand2 \comparator/C765  ( .a(\comparator/n1515 ), .b(\comparator/n1516 ), 
        .out(\comparator/N532 ) );
  nand2 \comparator/C766  ( .a(\comparator/n1517 ), .b(\comparator/n1518 ), 
        .out(\comparator/N530 ) );
  nand2 \comparator/C767  ( .a(\comparator/n1519 ), .b(\comparator/n1520 ), 
        .out(\comparator/N528 ) );
  nand2 \comparator/C768  ( .a(\comparator/n1521 ), .b(\comparator/n1522 ), 
        .out(\comparator/N526 ) );
  nand2 \comparator/C769  ( .a(\comparator/n1523 ), .b(\comparator/n1524 ), 
        .out(\comparator/N524 ) );
  nand2 \comparator/C770  ( .a(\comparator/n1525 ), .b(\comparator/n1526 ), 
        .out(\comparator/N522 ) );
  nand2 \comparator/C771  ( .a(\comparator/n1527 ), .b(\comparator/n1528 ), 
        .out(\comparator/N520 ) );
  nand2 \comparator/C772  ( .a(\comparator/n1529 ), .b(\comparator/n1530 ), 
        .out(\comparator/N518 ) );
  nand2 \comparator/C773  ( .a(\comparator/n1531 ), .b(\comparator/n1532 ), 
        .out(\comparator/N516 ) );
  nand2 \comparator/C774  ( .a(\comparator/n1533 ), .b(\comparator/n1534 ), 
        .out(\comparator/N514 ) );
  nand2 \comparator/C775  ( .a(\comparator/n1535 ), .b(\comparator/n1536 ), 
        .out(\comparator/N512 ) );
  nand2 \comparator/C776  ( .a(\comparator/n1537 ), .b(\comparator/n1538 ), 
        .out(\comparator/N510 ) );
  nand2 \comparator/C777  ( .a(\comparator/n1539 ), .b(\comparator/n1540 ), 
        .out(\comparator/N508 ) );
  nand2 \comparator/C778  ( .a(\comparator/n1541 ), .b(\comparator/n1542 ), 
        .out(\comparator/N506 ) );
  nand2 \comparator/C779  ( .a(\comparator/n1543 ), .b(\comparator/n1544 ), 
        .out(\comparator/N504 ) );
  nand2 \comparator/C780  ( .a(\comparator/n1545 ), .b(\comparator/n1546 ), 
        .out(\comparator/N502 ) );
  nand2 \comparator/C781  ( .a(\comparator/n1547 ), .b(\comparator/n1548 ), 
        .out(\comparator/N500 ) );
  nand2 \comparator/C782  ( .a(\comparator/n1549 ), .b(\comparator/n1550 ), 
        .out(\comparator/N498 ) );
  nand2 \comparator/C783  ( .a(\comparator/n1551 ), .b(\comparator/n1552 ), 
        .out(\comparator/N496 ) );
  nand2 \comparator/C784  ( .a(\comparator/n1553 ), .b(\comparator/n1554 ), 
        .out(\comparator/N494 ) );
  nand2 \comparator/C785  ( .a(\comparator/n1555 ), .b(\comparator/n1556 ), 
        .out(\comparator/N492 ) );
  nand2 \comparator/C786  ( .a(\comparator/n1557 ), .b(\comparator/n1558 ), 
        .out(\comparator/N490 ) );
  nand2 \comparator/C787  ( .a(\comparator/n1559 ), .b(\comparator/n1560 ), 
        .out(\comparator/N488 ) );
  nand2 \comparator/C788  ( .a(\comparator/n1561 ), .b(\comparator/n1562 ), 
        .out(\comparator/N486 ) );
  nand2 \comparator/C789  ( .a(\comparator/n1563 ), .b(\comparator/n1564 ), 
        .out(\comparator/N484 ) );
  nand2 \comparator/C790  ( .a(\comparator/n1565 ), .b(\comparator/n1566 ), 
        .out(\comparator/N482 ) );
  nand2 \comparator/C791  ( .a(\comparator/n1567 ), .b(\comparator/n1568 ), 
        .out(\comparator/N480 ) );
  nand2 \comparator/C792  ( .a(\comparator/n1569 ), .b(\comparator/n1570 ), 
        .out(\comparator/N478 ) );
  nand2 \comparator/C793  ( .a(\comparator/n1571 ), .b(\comparator/n1572 ), 
        .out(\comparator/N476 ) );
  nand2 \comparator/C794  ( .a(\comparator/n1573 ), .b(\comparator/n1574 ), 
        .out(\comparator/N474 ) );
  nand2 \comparator/C795  ( .a(\comparator/n1575 ), .b(\comparator/n1576 ), 
        .out(\comparator/N472 ) );
  nand2 \comparator/C796  ( .a(\comparator/n1577 ), .b(\comparator/n1578 ), 
        .out(\comparator/N470 ) );
  nand2 \comparator/C797  ( .a(\comparator/n1579 ), .b(\comparator/n1580 ), 
        .out(\comparator/N468 ) );
  nand2 \comparator/C798  ( .a(\comparator/n1581 ), .b(\comparator/n1582 ), 
        .out(\comparator/N466 ) );
  nand2 \comparator/C799  ( .a(\comparator/n1583 ), .b(\comparator/n1584 ), 
        .out(\comparator/N464 ) );
  nand2 \comparator/C800  ( .a(\comparator/n1585 ), .b(\comparator/n1586 ), 
        .out(\comparator/N462 ) );
  nand2 \comparator/C801  ( .a(\comparator/n1587 ), .b(\comparator/n1588 ), 
        .out(\comparator/N460 ) );
  nand2 \comparator/C802  ( .a(\comparator/n1589 ), .b(\comparator/n1590 ), 
        .out(\comparator/N458 ) );
  nand2 \comparator/C803  ( .a(\comparator/n1591 ), .b(\comparator/n1592 ), 
        .out(\comparator/N456 ) );
  nand2 \comparator/C804  ( .a(\comparator/n1593 ), .b(\comparator/n1594 ), 
        .out(\comparator/N454 ) );
  nand2 \comparator/C805  ( .a(\comparator/n1595 ), .b(\comparator/n1596 ), 
        .out(\comparator/N452 ) );
  nand2 \comparator/C806  ( .a(\comparator/n1597 ), .b(\comparator/n1598 ), 
        .out(\comparator/N450 ) );
  nand2 \comparator/C807  ( .a(\comparator/n1599 ), .b(\comparator/n1600 ), 
        .out(\comparator/N448 ) );
  nand2 \comparator/C808  ( .a(\comparator/n1601 ), .b(\comparator/n1602 ), 
        .out(\comparator/N446 ) );
  nand2 \comparator/C809  ( .a(\comparator/n1603 ), .b(\comparator/n1604 ), 
        .out(\comparator/N444 ) );
  nand2 \comparator/C810  ( .a(\comparator/n1605 ), .b(\comparator/n1606 ), 
        .out(\comparator/N442 ) );
  nand2 \comparator/C811  ( .a(\comparator/n1607 ), .b(\comparator/n1608 ), 
        .out(\comparator/N440 ) );
  nand2 \comparator/C812  ( .a(\comparator/n1609 ), .b(\comparator/n1610 ), 
        .out(\comparator/N438 ) );
  nand2 \comparator/C813  ( .a(\comparator/n1611 ), .b(\comparator/n1612 ), 
        .out(\comparator/N436 ) );
  nand2 \comparator/C814  ( .a(\comparator/n1613 ), .b(\comparator/n1614 ), 
        .out(\comparator/N434 ) );
  nand2 \comparator/C815  ( .a(\comparator/n1615 ), .b(\comparator/n1616 ), 
        .out(\comparator/N432 ) );
  nand2 \comparator/C816  ( .a(\comparator/n1617 ), .b(\comparator/n1618 ), 
        .out(\comparator/N430 ) );
  nand2 \comparator/C817  ( .a(\comparator/n1619 ), .b(\comparator/n1620 ), 
        .out(\comparator/N428 ) );
  nand2 \comparator/C818  ( .a(\comparator/n1621 ), .b(\comparator/n1622 ), 
        .out(\comparator/N426 ) );
  nand2 \comparator/C819  ( .a(\comparator/n1623 ), .b(\comparator/n1624 ), 
        .out(\comparator/N424 ) );
  nand2 \comparator/C820  ( .a(\comparator/n1625 ), .b(\comparator/n1626 ), 
        .out(\comparator/N422 ) );
  nand2 \comparator/C821  ( .a(\comparator/n1627 ), .b(\comparator/n1628 ), 
        .out(\comparator/N420 ) );
  nand2 \comparator/C822  ( .a(\comparator/n1629 ), .b(\comparator/n1630 ), 
        .out(\comparator/N418 ) );
  nand2 \comparator/C823  ( .a(\comparator/n1631 ), .b(\comparator/n1632 ), 
        .out(\comparator/N416 ) );
  nand2 \comparator/C824  ( .a(\comparator/n1633 ), .b(\comparator/n1634 ), 
        .out(\comparator/N414 ) );
  nand2 \comparator/C825  ( .a(\comparator/n1635 ), .b(\comparator/n1636 ), 
        .out(\comparator/N412 ) );
  nand2 \comparator/C826  ( .a(\comparator/n1637 ), .b(\comparator/n1638 ), 
        .out(\comparator/N410 ) );
  nand2 \comparator/C827  ( .a(\comparator/n1639 ), .b(\comparator/n1640 ), 
        .out(\comparator/N408 ) );
  nand2 \comparator/C828  ( .a(\comparator/n1641 ), .b(\comparator/n1642 ), 
        .out(\comparator/N406 ) );
  nand2 \comparator/C829  ( .a(\comparator/n1643 ), .b(\comparator/n1644 ), 
        .out(\comparator/N404 ) );
  nand2 \comparator/C830  ( .a(\comparator/n1645 ), .b(\comparator/n1646 ), 
        .out(\comparator/N402 ) );
  nand2 \comparator/C831  ( .a(\comparator/n1647 ), .b(\comparator/n1648 ), 
        .out(\comparator/N400 ) );
  nand2 \comparator/C832  ( .a(\comparator/n1649 ), .b(\comparator/n1650 ), 
        .out(\comparator/N398 ) );
  nand2 \comparator/C833  ( .a(\comparator/n1651 ), .b(\comparator/n1652 ), 
        .out(\comparator/N396 ) );
  nand2 \comparator/C834  ( .a(\comparator/n1653 ), .b(\comparator/n1654 ), 
        .out(\comparator/N394 ) );
  nand2 \comparator/C835  ( .a(\comparator/n1655 ), .b(\comparator/n1656 ), 
        .out(\comparator/N392 ) );
  nand2 \comparator/C836  ( .a(\comparator/n1657 ), .b(\comparator/n1658 ), 
        .out(\comparator/N390 ) );
  nand2 \comparator/C837  ( .a(\comparator/n1659 ), .b(\comparator/n1660 ), 
        .out(\comparator/N388 ) );
  nand2 \comparator/C838  ( .a(\comparator/n1661 ), .b(\comparator/n1662 ), 
        .out(\comparator/N386 ) );
  nand2 \comparator/C839  ( .a(\comparator/n1663 ), .b(\comparator/n1664 ), 
        .out(\comparator/N384 ) );
  nand2 \comparator/C840  ( .a(\comparator/n1665 ), .b(\comparator/n1666 ), 
        .out(\comparator/N382 ) );
  nand2 \comparator/C841  ( .a(\comparator/n1667 ), .b(\comparator/n1668 ), 
        .out(\comparator/N380 ) );
  nand2 \comparator/C842  ( .a(\comparator/n1669 ), .b(\comparator/n1670 ), 
        .out(\comparator/N378 ) );
  nand2 \comparator/C843  ( .a(\comparator/n1671 ), .b(\comparator/n1672 ), 
        .out(\comparator/N376 ) );
  nand2 \comparator/C844  ( .a(\comparator/n1673 ), .b(\comparator/n1674 ), 
        .out(\comparator/N374 ) );
  nand2 \comparator/C845  ( .a(\comparator/n1675 ), .b(\comparator/n1676 ), 
        .out(\comparator/N372 ) );
  nand2 \comparator/C846  ( .a(\comparator/n1677 ), .b(\comparator/n1678 ), 
        .out(\comparator/N370 ) );
  nand2 \comparator/C847  ( .a(\comparator/n1679 ), .b(\comparator/n1680 ), 
        .out(\comparator/N368 ) );
  nand2 \comparator/C848  ( .a(\comparator/n1681 ), .b(\comparator/n1682 ), 
        .out(\comparator/N366 ) );
  nand2 \comparator/C849  ( .a(\comparator/n1683 ), .b(\comparator/n1684 ), 
        .out(\comparator/N364 ) );
  nand2 \comparator/C850  ( .a(\comparator/n1685 ), .b(\comparator/n1686 ), 
        .out(\comparator/N362 ) );
  nand2 \comparator/C851  ( .a(\comparator/n1687 ), .b(\comparator/n1688 ), 
        .out(\comparator/N360 ) );
  nand2 \comparator/C852  ( .a(\comparator/n1689 ), .b(\comparator/n1690 ), 
        .out(\comparator/N358 ) );
  nand2 \comparator/C853  ( .a(\comparator/n1691 ), .b(\comparator/n1692 ), 
        .out(\comparator/N356 ) );
  nand2 \comparator/C854  ( .a(\comparator/n1693 ), .b(\comparator/n1694 ), 
        .out(\comparator/N354 ) );
  nand2 \comparator/C855  ( .a(\comparator/n1695 ), .b(\comparator/n1696 ), 
        .out(\comparator/N352 ) );
  nand2 \comparator/C856  ( .a(\comparator/n1697 ), .b(\comparator/n1698 ), 
        .out(\comparator/N350 ) );
  nand2 \comparator/C857  ( .a(\comparator/n1699 ), .b(\comparator/n1700 ), 
        .out(\comparator/N348 ) );
  nand2 \comparator/C858  ( .a(\comparator/n1701 ), .b(\comparator/n1702 ), 
        .out(\comparator/N346 ) );
  nand2 \comparator/C859  ( .a(\comparator/n1703 ), .b(\comparator/n1704 ), 
        .out(\comparator/N344 ) );
  nand2 \comparator/C860  ( .a(\comparator/n1705 ), .b(\comparator/n1706 ), 
        .out(\comparator/N342 ) );
  nand2 \comparator/C861  ( .a(\comparator/n1707 ), .b(\comparator/n1708 ), 
        .out(\comparator/N340 ) );
  nand2 \comparator/C862  ( .a(\comparator/n1709 ), .b(\comparator/n1710 ), 
        .out(\comparator/N338 ) );
  nand2 \comparator/C863  ( .a(\comparator/n1711 ), .b(\comparator/n1712 ), 
        .out(\comparator/N336 ) );
  nand2 \comparator/C864  ( .a(\comparator/n1713 ), .b(\comparator/n1714 ), 
        .out(\comparator/N334 ) );
  nand2 \comparator/C865  ( .a(\comparator/n1715 ), .b(\comparator/n1716 ), 
        .out(\comparator/N332 ) );
  nand2 \comparator/C866  ( .a(\comparator/n1717 ), .b(\comparator/n1718 ), 
        .out(\comparator/N330 ) );
  nand2 \comparator/C867  ( .a(\comparator/n1719 ), .b(\comparator/n1720 ), 
        .out(\comparator/N328 ) );
  nand2 \comparator/C868  ( .a(\comparator/n1721 ), .b(\comparator/n1722 ), 
        .out(\comparator/N326 ) );
  nand2 \comparator/C869  ( .a(\comparator/n1723 ), .b(\comparator/n1724 ), 
        .out(\comparator/N324 ) );
  nand2 \comparator/C870  ( .a(\comparator/n1725 ), .b(\comparator/n1726 ), 
        .out(\comparator/N322 ) );
  nand2 \comparator/C871  ( .a(\comparator/n1727 ), .b(\comparator/n1728 ), 
        .out(\comparator/N320 ) );
  nand2 \comparator/C872  ( .a(\comparator/n1729 ), .b(\comparator/n1730 ), 
        .out(\comparator/N318 ) );
  nand2 \comparator/C873  ( .a(\comparator/n1731 ), .b(\comparator/n1732 ), 
        .out(\comparator/N316 ) );
  nand2 \comparator/C874  ( .a(\comparator/n1733 ), .b(\comparator/n1734 ), 
        .out(\comparator/N314 ) );
  nand2 \comparator/C875  ( .a(\comparator/n1735 ), .b(\comparator/n1736 ), 
        .out(\comparator/N312 ) );
  nand2 \comparator/C876  ( .a(\comparator/n1737 ), .b(\comparator/n1738 ), 
        .out(\comparator/N310 ) );
  nand2 \comparator/C877  ( .a(\comparator/n1739 ), .b(\comparator/n1740 ), 
        .out(\comparator/N308 ) );
  nand2 \comparator/C878  ( .a(\comparator/n1741 ), .b(\comparator/n1742 ), 
        .out(\comparator/N306 ) );
  nand2 \comparator/C879  ( .a(\comparator/n1743 ), .b(\comparator/n1744 ), 
        .out(\comparator/N304 ) );
  nand2 \comparator/C880  ( .a(\comparator/n1745 ), .b(\comparator/n1746 ), 
        .out(\comparator/N302 ) );
  nand2 \comparator/C881  ( .a(\comparator/n1747 ), .b(\comparator/n1748 ), 
        .out(\comparator/N300 ) );
  nand2 \comparator/C882  ( .a(\comparator/n1749 ), .b(\comparator/n1750 ), 
        .out(\comparator/N298 ) );
  nand2 \comparator/C883  ( .a(\comparator/n1751 ), .b(\comparator/n1752 ), 
        .out(\comparator/N296 ) );
  nand2 \comparator/C884  ( .a(\comparator/n1753 ), .b(\comparator/n1754 ), 
        .out(\comparator/N294 ) );
  nand2 \comparator/C885  ( .a(\comparator/n1755 ), .b(\comparator/n1756 ), 
        .out(\comparator/N292 ) );
  nand2 \comparator/C886  ( .a(\comparator/n1757 ), .b(\comparator/n1758 ), 
        .out(\comparator/N290 ) );
  nand2 \comparator/C887  ( .a(\comparator/n1759 ), .b(\comparator/n1760 ), 
        .out(\comparator/N288 ) );
  nand2 \comparator/C888  ( .a(\comparator/n1761 ), .b(\comparator/n1762 ), 
        .out(\comparator/N286 ) );
  nand2 \comparator/C889  ( .a(\comparator/n1763 ), .b(\comparator/n1764 ), 
        .out(\comparator/N284 ) );
  nand2 \comparator/C890  ( .a(\comparator/n1765 ), .b(\comparator/n1766 ), 
        .out(\comparator/N282 ) );
  nand2 \comparator/C891  ( .a(\comparator/n1767 ), .b(\comparator/n1768 ), 
        .out(\comparator/N280 ) );
  nand2 \comparator/C892  ( .a(\comparator/n1769 ), .b(\comparator/n1770 ), 
        .out(\comparator/N278 ) );
  nand2 \comparator/C893  ( .a(\comparator/n1771 ), .b(\comparator/n1772 ), 
        .out(\comparator/N276 ) );
  nand2 \comparator/C894  ( .a(\comparator/n1773 ), .b(\comparator/n1774 ), 
        .out(\comparator/N274 ) );
  nand2 \comparator/C895  ( .a(\comparator/n1775 ), .b(\comparator/n1776 ), 
        .out(\comparator/N272 ) );
  nand2 \comparator/C896  ( .a(\comparator/n1777 ), .b(\comparator/n1778 ), 
        .out(\comparator/N270 ) );
  nand2 \comparator/C897  ( .a(\comparator/n1779 ), .b(\comparator/n1780 ), 
        .out(\comparator/N268 ) );
  nand2 \comparator/C898  ( .a(\comparator/n1781 ), .b(\comparator/n1782 ), 
        .out(\comparator/N266 ) );
  nand2 \comparator/C899  ( .a(\comparator/n1783 ), .b(\comparator/n1784 ), 
        .out(\comparator/N264 ) );
  nand2 \comparator/C900  ( .a(\comparator/n1785 ), .b(\comparator/n1786 ), 
        .out(\comparator/N262 ) );
  nand2 \comparator/C901  ( .a(\comparator/n1787 ), .b(\comparator/n1788 ), 
        .out(\comparator/N260 ) );
  nand2 \comparator/C902  ( .a(\comparator/n1789 ), .b(\comparator/n1790 ), 
        .out(\comparator/N258 ) );
  nand2 \comparator/C903  ( .a(\comparator/n1791 ), .b(\comparator/n1792 ), 
        .out(\comparator/N256 ) );
  nand2 \comparator/C904  ( .a(\comparator/n1793 ), .b(\comparator/n1794 ), 
        .out(\comparator/N254 ) );
  nand2 \comparator/C905  ( .a(\comparator/n1795 ), .b(\comparator/n1796 ), 
        .out(\comparator/N252 ) );
  nand2 \comparator/C906  ( .a(\comparator/n1797 ), .b(\comparator/n1798 ), 
        .out(\comparator/N250 ) );
  nand2 \comparator/C907  ( .a(\comparator/n1799 ), .b(\comparator/n1800 ), 
        .out(\comparator/N248 ) );
  nand2 \comparator/C908  ( .a(\comparator/n1801 ), .b(\comparator/n1802 ), 
        .out(\comparator/N246 ) );
  nand2 \comparator/C909  ( .a(\comparator/n1803 ), .b(\comparator/n1804 ), 
        .out(\comparator/N244 ) );
  nand2 \comparator/C910  ( .a(\comparator/n1805 ), .b(\comparator/n1806 ), 
        .out(\comparator/N242 ) );
  nand2 \comparator/C911  ( .a(\comparator/n1807 ), .b(\comparator/n1808 ), 
        .out(\comparator/N240 ) );
  nand2 \comparator/C912  ( .a(\comparator/n1809 ), .b(\comparator/n1810 ), 
        .out(\comparator/N238 ) );
  nand2 \comparator/C913  ( .a(\comparator/n1811 ), .b(\comparator/n1812 ), 
        .out(\comparator/N236 ) );
  nand2 \comparator/C914  ( .a(\comparator/n1813 ), .b(\comparator/n1814 ), 
        .out(\comparator/N234 ) );
  nand2 \comparator/C915  ( .a(\comparator/n1815 ), .b(\comparator/n1816 ), 
        .out(\comparator/N232 ) );
  nand2 \comparator/C916  ( .a(\comparator/n1817 ), .b(\comparator/n1818 ), 
        .out(\comparator/N230 ) );
  nand2 \comparator/C917  ( .a(\comparator/n1819 ), .b(\comparator/n1820 ), 
        .out(\comparator/N228 ) );
  nand2 \comparator/C918  ( .a(\comparator/n1821 ), .b(\comparator/n1822 ), 
        .out(\comparator/N226 ) );
  nand2 \comparator/C919  ( .a(\comparator/n1823 ), .b(\comparator/n1824 ), 
        .out(\comparator/N224 ) );
  nand2 \comparator/C920  ( .a(\comparator/n1825 ), .b(\comparator/n1826 ), 
        .out(\comparator/N222 ) );
  nand2 \comparator/C921  ( .a(\comparator/n1827 ), .b(\comparator/n1828 ), 
        .out(\comparator/N220 ) );
  nand2 \comparator/C922  ( .a(\comparator/n1829 ), .b(\comparator/n1830 ), 
        .out(\comparator/N218 ) );
  nand2 \comparator/C923  ( .a(\comparator/n1831 ), .b(\comparator/n1832 ), 
        .out(\comparator/N216 ) );
  nand2 \comparator/C924  ( .a(\comparator/n1833 ), .b(\comparator/n1834 ), 
        .out(\comparator/N214 ) );
  nand2 \comparator/C925  ( .a(\comparator/n1835 ), .b(\comparator/n1836 ), 
        .out(\comparator/N212 ) );
  nand2 \comparator/C926  ( .a(\comparator/n1837 ), .b(\comparator/n1838 ), 
        .out(\comparator/N210 ) );
  nand2 \comparator/C927  ( .a(\comparator/n1839 ), .b(\comparator/n1840 ), 
        .out(\comparator/N208 ) );
  nand2 \comparator/C928  ( .a(\comparator/n1841 ), .b(\comparator/n1842 ), 
        .out(\comparator/N206 ) );
  nand2 \comparator/C929  ( .a(\comparator/n1843 ), .b(\comparator/n1844 ), 
        .out(\comparator/N204 ) );
  nand2 \comparator/C930  ( .a(\comparator/n1845 ), .b(\comparator/n1846 ), 
        .out(\comparator/N202 ) );
  nand2 \comparator/C931  ( .a(\comparator/n1847 ), .b(\comparator/n1848 ), 
        .out(\comparator/N200 ) );
  nand2 \comparator/C932  ( .a(\comparator/n1849 ), .b(\comparator/n1850 ), 
        .out(\comparator/N198 ) );
  nand2 \comparator/C933  ( .a(\comparator/n1851 ), .b(\comparator/n1852 ), 
        .out(\comparator/N196 ) );
  nand2 \comparator/C934  ( .a(\comparator/n1853 ), .b(\comparator/n1854 ), 
        .out(\comparator/N194 ) );
  nand2 \comparator/C935  ( .a(\comparator/n1855 ), .b(\comparator/n1856 ), 
        .out(\comparator/N192 ) );
  nand2 \comparator/C936  ( .a(\comparator/n1857 ), .b(\comparator/n1858 ), 
        .out(\comparator/N190 ) );
  nand2 \comparator/C937  ( .a(\comparator/n1859 ), .b(\comparator/n1860 ), 
        .out(\comparator/N188 ) );
  nand2 \comparator/C938  ( .a(\comparator/n1861 ), .b(\comparator/n1862 ), 
        .out(\comparator/N186 ) );
  nand2 \comparator/C939  ( .a(\comparator/n1863 ), .b(\comparator/n1864 ), 
        .out(\comparator/N184 ) );
  nand2 \comparator/C940  ( .a(\comparator/n1865 ), .b(\comparator/n1866 ), 
        .out(\comparator/N182 ) );
  nand2 \comparator/C941  ( .a(\comparator/n1867 ), .b(\comparator/n1868 ), 
        .out(\comparator/N180 ) );
  nand2 \comparator/C942  ( .a(\comparator/n1869 ), .b(\comparator/n1870 ), 
        .out(\comparator/N178 ) );
  nand2 \comparator/C943  ( .a(\comparator/n1871 ), .b(\comparator/n1872 ), 
        .out(\comparator/N176 ) );
  nand2 \comparator/C944  ( .a(\comparator/n1873 ), .b(\comparator/n1874 ), 
        .out(\comparator/N174 ) );
  nand2 \comparator/C945  ( .a(\comparator/n1875 ), .b(\comparator/n1876 ), 
        .out(\comparator/N172 ) );
  nand2 \comparator/C946  ( .a(\comparator/n1877 ), .b(\comparator/n1878 ), 
        .out(\comparator/N170 ) );
  nand2 \comparator/C947  ( .a(\comparator/n1879 ), .b(\comparator/n1880 ), 
        .out(\comparator/N168 ) );
  nand2 \comparator/C948  ( .a(\comparator/n1881 ), .b(\comparator/n1882 ), 
        .out(\comparator/N166 ) );
  nand2 \comparator/C949  ( .a(\comparator/n1883 ), .b(\comparator/n1884 ), 
        .out(\comparator/N164 ) );
  nand2 \comparator/C950  ( .a(\comparator/n1885 ), .b(\comparator/n1886 ), 
        .out(\comparator/N162 ) );
  nand2 \comparator/C951  ( .a(\comparator/n1887 ), .b(\comparator/n1888 ), 
        .out(\comparator/N160 ) );
  nand2 \comparator/C952  ( .a(\comparator/n1889 ), .b(\comparator/n1890 ), 
        .out(\comparator/N158 ) );
  nand2 \comparator/C953  ( .a(\comparator/n1891 ), .b(\comparator/n1892 ), 
        .out(\comparator/N156 ) );
  nand2 \comparator/C954  ( .a(\comparator/n1893 ), .b(\comparator/n1894 ), 
        .out(\comparator/N154 ) );
  nand2 \comparator/C955  ( .a(\comparator/n1895 ), .b(\comparator/n1896 ), 
        .out(\comparator/N152 ) );
  nand2 \comparator/C956  ( .a(\comparator/n1897 ), .b(\comparator/n1898 ), 
        .out(\comparator/N150 ) );
  nand2 \comparator/C957  ( .a(\comparator/n1899 ), .b(\comparator/n1900 ), 
        .out(\comparator/N148 ) );
  nand2 \comparator/C958  ( .a(\comparator/n1901 ), .b(\comparator/n1902 ), 
        .out(\comparator/N146 ) );
  nand2 \comparator/C959  ( .a(\comparator/n1903 ), .b(\comparator/n1904 ), 
        .out(\comparator/N144 ) );
  nand2 \comparator/C960  ( .a(\comparator/n1905 ), .b(\comparator/n1906 ), 
        .out(\comparator/N142 ) );
  nand2 \comparator/C961  ( .a(\comparator/n1907 ), .b(\comparator/n1908 ), 
        .out(\comparator/N140 ) );
  nand2 \comparator/C962  ( .a(\comparator/n1909 ), .b(\comparator/n1910 ), 
        .out(\comparator/N138 ) );
  nand2 \comparator/C963  ( .a(\comparator/n1911 ), .b(\comparator/n1912 ), 
        .out(\comparator/N136 ) );
  nand2 \comparator/C964  ( .a(\comparator/n1913 ), .b(\comparator/n1914 ), 
        .out(\comparator/N134 ) );
  nand2 \comparator/C965  ( .a(\comparator/n1915 ), .b(\comparator/n1916 ), 
        .out(\comparator/N132 ) );
  nand2 \comparator/C966  ( .a(\comparator/n1917 ), .b(\comparator/n1918 ), 
        .out(\comparator/N130 ) );
  nand2 \comparator/C967  ( .a(\comparator/n1919 ), .b(\comparator/n1920 ), 
        .out(\comparator/N128 ) );
  nand2 \comparator/C968  ( .a(\comparator/n1921 ), .b(\comparator/n1922 ), 
        .out(\comparator/N126 ) );
  nand2 \comparator/C969  ( .a(\comparator/n1923 ), .b(\comparator/n1924 ), 
        .out(\comparator/N124 ) );
  nand2 \comparator/C970  ( .a(\comparator/n1925 ), .b(\comparator/n1926 ), 
        .out(\comparator/N122 ) );
  nand2 \comparator/C971  ( .a(\comparator/n1927 ), .b(\comparator/n1928 ), 
        .out(\comparator/N120 ) );
  nand2 \comparator/C972  ( .a(\comparator/n1929 ), .b(\comparator/n1930 ), 
        .out(\comparator/N118 ) );
  nand2 \comparator/C973  ( .a(\comparator/n1931 ), .b(\comparator/n1932 ), 
        .out(\comparator/N116 ) );
  nand2 \comparator/C974  ( .a(\comparator/n1933 ), .b(\comparator/n1934 ), 
        .out(\comparator/N114 ) );
  nand2 \comparator/C975  ( .a(\comparator/n1935 ), .b(\comparator/n1936 ), 
        .out(\comparator/N112 ) );
  nand2 \comparator/C976  ( .a(\comparator/n1937 ), .b(\comparator/n1938 ), 
        .out(\comparator/N110 ) );
  nand2 \comparator/C977  ( .a(\comparator/n1939 ), .b(\comparator/n1940 ), 
        .out(\comparator/N108 ) );
  nand2 \comparator/C978  ( .a(\comparator/n1941 ), .b(\comparator/n1942 ), 
        .out(\comparator/N106 ) );
  nand2 \comparator/C979  ( .a(\comparator/n1943 ), .b(\comparator/n1944 ), 
        .out(\comparator/N104 ) );
  nand2 \comparator/C980  ( .a(\comparator/n1945 ), .b(\comparator/n1946 ), 
        .out(\comparator/N102 ) );
  nand2 \comparator/C981  ( .a(\comparator/n1947 ), .b(\comparator/n1948 ), 
        .out(\comparator/N100 ) );
  nand2 \comparator/C982  ( .a(\comparator/n1949 ), .b(\comparator/n1950 ), 
        .out(\comparator/N98 ) );
  nand2 \comparator/C983  ( .a(\comparator/n1951 ), .b(\comparator/n1952 ), 
        .out(\comparator/N96 ) );
  nand2 \comparator/C984  ( .a(\comparator/n1953 ), .b(\comparator/n1954 ), 
        .out(\comparator/N94 ) );
  nand2 \comparator/C985  ( .a(\comparator/n1955 ), .b(\comparator/n1956 ), 
        .out(\comparator/N92 ) );
  nand2 \comparator/C986  ( .a(\comparator/n1957 ), .b(\comparator/n1958 ), 
        .out(\comparator/N90 ) );
  nand2 \comparator/C987  ( .a(\comparator/n1959 ), .b(\comparator/n1960 ), 
        .out(\comparator/N88 ) );
  nand2 \comparator/C988  ( .a(\comparator/n1961 ), .b(\comparator/n1962 ), 
        .out(\comparator/N86 ) );
  nand2 \comparator/C989  ( .a(\comparator/n1963 ), .b(\comparator/n1964 ), 
        .out(\comparator/N84 ) );
  nand2 \comparator/C990  ( .a(\comparator/n1965 ), .b(\comparator/n1966 ), 
        .out(\comparator/N82 ) );
  nand2 \comparator/C991  ( .a(\comparator/n1967 ), .b(\comparator/n1968 ), 
        .out(\comparator/N80 ) );
  nand2 \comparator/C992  ( .a(\comparator/n1969 ), .b(\comparator/n1970 ), 
        .out(\comparator/N78 ) );
  nand2 \comparator/C993  ( .a(\comparator/n1971 ), .b(\comparator/n1972 ), 
        .out(\comparator/N76 ) );
  nand2 \comparator/C994  ( .a(\comparator/n1973 ), .b(\comparator/n1974 ), 
        .out(\comparator/N74 ) );
  nand2 \comparator/C995  ( .a(\comparator/n1975 ), .b(\comparator/n1976 ), 
        .out(\comparator/N72 ) );
  nand2 \comparator/C996  ( .a(\comparator/n1977 ), .b(\comparator/n1978 ), 
        .out(\comparator/N70 ) );
  nand2 \comparator/C997  ( .a(\comparator/n1979 ), .b(\comparator/n1980 ), 
        .out(\comparator/N68 ) );
  nand2 \comparator/C998  ( .a(\comparator/n1981 ), .b(\comparator/n1982 ), 
        .out(\comparator/N66 ) );
  nand2 \comparator/C999  ( .a(\comparator/n1983 ), .b(\comparator/n1984 ), 
        .out(\comparator/N64 ) );
  nand2 \comparator/C1000  ( .a(\comparator/n1985 ), .b(\comparator/n1986 ), 
        .out(\comparator/N62 ) );
  nand2 \comparator/C1001  ( .a(\comparator/n1987 ), .b(\comparator/n1988 ), 
        .out(\comparator/N60 ) );
  nand2 \comparator/C1002  ( .a(\comparator/n1989 ), .b(\comparator/n1990 ), 
        .out(\comparator/N58 ) );
  nand2 \comparator/C1003  ( .a(\comparator/n1991 ), .b(\comparator/n1992 ), 
        .out(\comparator/N56 ) );
  nand2 \comparator/C1004  ( .a(\comparator/n1993 ), .b(\comparator/n1994 ), 
        .out(\comparator/N54 ) );
  nand2 \comparator/C1005  ( .a(\comparator/n1995 ), .b(\comparator/n1996 ), 
        .out(\comparator/N52 ) );
  nand2 \comparator/C1006  ( .a(\comparator/n1997 ), .b(\comparator/n1998 ), 
        .out(\comparator/N50 ) );
  nand2 \comparator/C1007  ( .a(\comparator/n1999 ), .b(\comparator/n2000 ), 
        .out(\comparator/N48 ) );
  nand2 \comparator/C1008  ( .a(\comparator/n2001 ), .b(\comparator/n2002 ), 
        .out(\comparator/N46 ) );
  nand2 \comparator/C1009  ( .a(\comparator/n2003 ), .b(\comparator/n2004 ), 
        .out(\comparator/N44 ) );
  nand2 \comparator/C1010  ( .a(\comparator/n2005 ), .b(\comparator/n2006 ), 
        .out(\comparator/N42 ) );
  nand2 \comparator/C1011  ( .a(\comparator/n2007 ), .b(\comparator/n2008 ), 
        .out(\comparator/N40 ) );
  nand2 \comparator/C1012  ( .a(\comparator/n2009 ), .b(\comparator/n2010 ), 
        .out(\comparator/N38 ) );
  nand2 \comparator/C1013  ( .a(\comparator/n2011 ), .b(\comparator/n2012 ), 
        .out(\comparator/N36 ) );
  nand2 \comparator/C1014  ( .a(\comparator/n2013 ), .b(\comparator/n2014 ), 
        .out(\comparator/N34 ) );
  nand2 \comparator/C1015  ( .a(\comparator/n2015 ), .b(\comparator/n2016 ), 
        .out(\comparator/N32 ) );
  nand2 \comparator/C1016  ( .a(\comparator/n2017 ), .b(\comparator/n2018 ), 
        .out(\comparator/N30 ) );
  nand2 \comparator/C1017  ( .a(\comparator/n2019 ), .b(\comparator/n2020 ), 
        .out(\comparator/N28 ) );
  nand2 \comparator/C1018  ( .a(\comparator/n2021 ), .b(\comparator/n2022 ), 
        .out(\comparator/N26 ) );
  nand2 \comparator/C1019  ( .a(\comparator/n2023 ), .b(\comparator/n2024 ), 
        .out(\comparator/N24 ) );
  nand2 \comparator/C1020  ( .a(\comparator/n2025 ), .b(\comparator/n2026 ), 
        .out(\comparator/N22 ) );
  nand2 \comparator/C1021  ( .a(\comparator/n2027 ), .b(\comparator/n2028 ), 
        .out(\comparator/N20 ) );
  nand2 \comparator/C1022  ( .a(\comparator/n2029 ), .b(\comparator/n2030 ), 
        .out(\comparator/N18 ) );
  nand2 \comparator/C1023  ( .a(\comparator/n2031 ), .b(\comparator/n2032 ), 
        .out(\comparator/N16 ) );
  nand2 \comparator/C1024  ( .a(\comparator/n2033 ), .b(\comparator/n2034 ), 
        .out(\comparator/N14 ) );
  nand2 \comparator/C1025  ( .a(\comparator/n2035 ), .b(\comparator/n2036 ), 
        .out(\comparator/N12 ) );
  nand2 \comparator/C1026  ( .a(\comparator/n2037 ), .b(\comparator/n2038 ), 
        .out(\comparator/N10 ) );
  nand2 \comparator/C1027  ( .a(\comparator/n2039 ), .b(\comparator/n2040 ), 
        .out(\comparator/N8 ) );
  nand2 \comparator/C1028  ( .a(\comparator/n2041 ), .b(\comparator/n2042 ), 
        .out(\comparator/N6 ) );
  nand2 \comparator/C1029  ( .a(\comparator/n2043 ), .b(\comparator/n2044 ), 
        .out(\comparator/N4 ) );
  nand2 \comparator/C1030  ( .a(\comparator/n2045 ), .b(\comparator/n2046 ), 
        .out(\comparator/N2 ) );
  xor2 \comparator/C1031  ( .a(a[1023]), .b(b[1023]), .out(\comparator/N0 ) );
  xor2 \comparator/C1032  ( .a(a[1022]), .b(b[1022]), .out(\comparator/N1 ) );
  xor2 \comparator/C1033  ( .a(a[1021]), .b(b[1021]), .out(\comparator/N3 ) );
  xor2 \comparator/C1034  ( .a(a[1020]), .b(b[1020]), .out(\comparator/N5 ) );
  xor2 \comparator/C1035  ( .a(a[1019]), .b(b[1019]), .out(\comparator/N7 ) );
  xor2 \comparator/C1036  ( .a(a[1018]), .b(b[1018]), .out(\comparator/N9 ) );
  xor2 \comparator/C1037  ( .a(a[1017]), .b(b[1017]), .out(\comparator/N11 )
         );
  xor2 \comparator/C1038  ( .a(a[1016]), .b(b[1016]), .out(\comparator/N13 )
         );
  xor2 \comparator/C1039  ( .a(a[1015]), .b(b[1015]), .out(\comparator/N15 )
         );
  xor2 \comparator/C1040  ( .a(a[1014]), .b(b[1014]), .out(\comparator/N17 )
         );
  xor2 \comparator/C1041  ( .a(a[1013]), .b(b[1013]), .out(\comparator/N19 )
         );
  xor2 \comparator/C1042  ( .a(a[1012]), .b(b[1012]), .out(\comparator/N21 )
         );
  xor2 \comparator/C1043  ( .a(a[1011]), .b(b[1011]), .out(\comparator/N23 )
         );
  xor2 \comparator/C1044  ( .a(a[1010]), .b(b[1010]), .out(\comparator/N25 )
         );
  xor2 \comparator/C1045  ( .a(a[1009]), .b(b[1009]), .out(\comparator/N27 )
         );
  xor2 \comparator/C1046  ( .a(a[1008]), .b(b[1008]), .out(\comparator/N29 )
         );
  xor2 \comparator/C1047  ( .a(a[1007]), .b(b[1007]), .out(\comparator/N31 )
         );
  xor2 \comparator/C1048  ( .a(a[1006]), .b(b[1006]), .out(\comparator/N33 )
         );
  xor2 \comparator/C1049  ( .a(a[1005]), .b(b[1005]), .out(\comparator/N35 )
         );
  xor2 \comparator/C1050  ( .a(a[1004]), .b(b[1004]), .out(\comparator/N37 )
         );
  xor2 \comparator/C1051  ( .a(a[1003]), .b(b[1003]), .out(\comparator/N39 )
         );
  xor2 \comparator/C1052  ( .a(a[1002]), .b(b[1002]), .out(\comparator/N41 )
         );
  xor2 \comparator/C1053  ( .a(a[1001]), .b(b[1001]), .out(\comparator/N43 )
         );
  xor2 \comparator/C1054  ( .a(a[1000]), .b(b[1000]), .out(\comparator/N45 )
         );
  xor2 \comparator/C1055  ( .a(a[999]), .b(b[999]), .out(\comparator/N47 ) );
  xor2 \comparator/C1056  ( .a(a[998]), .b(b[998]), .out(\comparator/N49 ) );
  xor2 \comparator/C1057  ( .a(a[997]), .b(b[997]), .out(\comparator/N51 ) );
  xor2 \comparator/C1058  ( .a(a[996]), .b(b[996]), .out(\comparator/N53 ) );
  xor2 \comparator/C1059  ( .a(a[995]), .b(b[995]), .out(\comparator/N55 ) );
  xor2 \comparator/C1060  ( .a(a[994]), .b(b[994]), .out(\comparator/N57 ) );
  xor2 \comparator/C1061  ( .a(a[993]), .b(b[993]), .out(\comparator/N59 ) );
  xor2 \comparator/C1062  ( .a(a[992]), .b(b[992]), .out(\comparator/N61 ) );
  xor2 \comparator/C1063  ( .a(a[991]), .b(b[991]), .out(\comparator/N63 ) );
  xor2 \comparator/C1064  ( .a(a[990]), .b(b[990]), .out(\comparator/N65 ) );
  xor2 \comparator/C1065  ( .a(a[989]), .b(b[989]), .out(\comparator/N67 ) );
  xor2 \comparator/C1066  ( .a(a[988]), .b(b[988]), .out(\comparator/N69 ) );
  xor2 \comparator/C1067  ( .a(a[987]), .b(b[987]), .out(\comparator/N71 ) );
  xor2 \comparator/C1068  ( .a(a[986]), .b(b[986]), .out(\comparator/N73 ) );
  xor2 \comparator/C1069  ( .a(a[985]), .b(b[985]), .out(\comparator/N75 ) );
  xor2 \comparator/C1070  ( .a(a[984]), .b(b[984]), .out(\comparator/N77 ) );
  xor2 \comparator/C1071  ( .a(a[983]), .b(b[983]), .out(\comparator/N79 ) );
  xor2 \comparator/C1072  ( .a(a[982]), .b(b[982]), .out(\comparator/N81 ) );
  xor2 \comparator/C1073  ( .a(a[981]), .b(b[981]), .out(\comparator/N83 ) );
  xor2 \comparator/C1074  ( .a(a[980]), .b(b[980]), .out(\comparator/N85 ) );
  xor2 \comparator/C1075  ( .a(a[979]), .b(b[979]), .out(\comparator/N87 ) );
  xor2 \comparator/C1076  ( .a(a[978]), .b(b[978]), .out(\comparator/N89 ) );
  xor2 \comparator/C1077  ( .a(a[977]), .b(b[977]), .out(\comparator/N91 ) );
  xor2 \comparator/C1078  ( .a(a[976]), .b(b[976]), .out(\comparator/N93 ) );
  xor2 \comparator/C1079  ( .a(a[975]), .b(b[975]), .out(\comparator/N95 ) );
  xor2 \comparator/C1080  ( .a(a[974]), .b(b[974]), .out(\comparator/N97 ) );
  xor2 \comparator/C1081  ( .a(a[973]), .b(b[973]), .out(\comparator/N99 ) );
  xor2 \comparator/C1082  ( .a(a[972]), .b(b[972]), .out(\comparator/N101 ) );
  xor2 \comparator/C1083  ( .a(a[971]), .b(b[971]), .out(\comparator/N103 ) );
  xor2 \comparator/C1084  ( .a(a[970]), .b(b[970]), .out(\comparator/N105 ) );
  xor2 \comparator/C1085  ( .a(a[969]), .b(b[969]), .out(\comparator/N107 ) );
  xor2 \comparator/C1086  ( .a(a[968]), .b(b[968]), .out(\comparator/N109 ) );
  xor2 \comparator/C1087  ( .a(a[967]), .b(b[967]), .out(\comparator/N111 ) );
  xor2 \comparator/C1088  ( .a(a[966]), .b(b[966]), .out(\comparator/N113 ) );
  xor2 \comparator/C1089  ( .a(a[965]), .b(b[965]), .out(\comparator/N115 ) );
  xor2 \comparator/C1090  ( .a(a[964]), .b(b[964]), .out(\comparator/N117 ) );
  xor2 \comparator/C1091  ( .a(a[963]), .b(b[963]), .out(\comparator/N119 ) );
  xor2 \comparator/C1092  ( .a(a[962]), .b(b[962]), .out(\comparator/N121 ) );
  xor2 \comparator/C1093  ( .a(a[961]), .b(b[961]), .out(\comparator/N123 ) );
  xor2 \comparator/C1094  ( .a(a[960]), .b(b[960]), .out(\comparator/N125 ) );
  xor2 \comparator/C1095  ( .a(a[959]), .b(b[959]), .out(\comparator/N127 ) );
  xor2 \comparator/C1096  ( .a(a[958]), .b(b[958]), .out(\comparator/N129 ) );
  xor2 \comparator/C1097  ( .a(a[957]), .b(b[957]), .out(\comparator/N131 ) );
  xor2 \comparator/C1098  ( .a(a[956]), .b(b[956]), .out(\comparator/N133 ) );
  xor2 \comparator/C1099  ( .a(a[955]), .b(b[955]), .out(\comparator/N135 ) );
  xor2 \comparator/C1100  ( .a(a[954]), .b(b[954]), .out(\comparator/N137 ) );
  xor2 \comparator/C1101  ( .a(a[953]), .b(b[953]), .out(\comparator/N139 ) );
  xor2 \comparator/C1102  ( .a(a[952]), .b(b[952]), .out(\comparator/N141 ) );
  xor2 \comparator/C1103  ( .a(a[951]), .b(b[951]), .out(\comparator/N143 ) );
  xor2 \comparator/C1104  ( .a(a[950]), .b(b[950]), .out(\comparator/N145 ) );
  xor2 \comparator/C1105  ( .a(a[949]), .b(b[949]), .out(\comparator/N147 ) );
  xor2 \comparator/C1106  ( .a(a[948]), .b(b[948]), .out(\comparator/N149 ) );
  xor2 \comparator/C1107  ( .a(a[947]), .b(b[947]), .out(\comparator/N151 ) );
  xor2 \comparator/C1108  ( .a(a[946]), .b(b[946]), .out(\comparator/N153 ) );
  xor2 \comparator/C1109  ( .a(a[945]), .b(b[945]), .out(\comparator/N155 ) );
  xor2 \comparator/C1110  ( .a(a[944]), .b(b[944]), .out(\comparator/N157 ) );
  xor2 \comparator/C1111  ( .a(a[943]), .b(b[943]), .out(\comparator/N159 ) );
  xor2 \comparator/C1112  ( .a(a[942]), .b(b[942]), .out(\comparator/N161 ) );
  xor2 \comparator/C1113  ( .a(a[941]), .b(b[941]), .out(\comparator/N163 ) );
  xor2 \comparator/C1114  ( .a(a[940]), .b(b[940]), .out(\comparator/N165 ) );
  xor2 \comparator/C1115  ( .a(a[939]), .b(b[939]), .out(\comparator/N167 ) );
  xor2 \comparator/C1116  ( .a(a[938]), .b(b[938]), .out(\comparator/N169 ) );
  xor2 \comparator/C1117  ( .a(a[937]), .b(b[937]), .out(\comparator/N171 ) );
  xor2 \comparator/C1118  ( .a(a[936]), .b(b[936]), .out(\comparator/N173 ) );
  xor2 \comparator/C1119  ( .a(a[935]), .b(b[935]), .out(\comparator/N175 ) );
  xor2 \comparator/C1120  ( .a(a[934]), .b(b[934]), .out(\comparator/N177 ) );
  xor2 \comparator/C1121  ( .a(a[933]), .b(b[933]), .out(\comparator/N179 ) );
  xor2 \comparator/C1122  ( .a(a[932]), .b(b[932]), .out(\comparator/N181 ) );
  xor2 \comparator/C1123  ( .a(a[931]), .b(b[931]), .out(\comparator/N183 ) );
  xor2 \comparator/C1124  ( .a(a[930]), .b(b[930]), .out(\comparator/N185 ) );
  xor2 \comparator/C1125  ( .a(a[929]), .b(b[929]), .out(\comparator/N187 ) );
  xor2 \comparator/C1126  ( .a(a[928]), .b(b[928]), .out(\comparator/N189 ) );
  xor2 \comparator/C1127  ( .a(a[927]), .b(b[927]), .out(\comparator/N191 ) );
  xor2 \comparator/C1128  ( .a(a[926]), .b(b[926]), .out(\comparator/N193 ) );
  xor2 \comparator/C1129  ( .a(a[925]), .b(b[925]), .out(\comparator/N195 ) );
  xor2 \comparator/C1130  ( .a(a[924]), .b(b[924]), .out(\comparator/N197 ) );
  xor2 \comparator/C1131  ( .a(a[923]), .b(b[923]), .out(\comparator/N199 ) );
  xor2 \comparator/C1132  ( .a(a[922]), .b(b[922]), .out(\comparator/N201 ) );
  xor2 \comparator/C1133  ( .a(a[921]), .b(b[921]), .out(\comparator/N203 ) );
  xor2 \comparator/C1134  ( .a(a[920]), .b(b[920]), .out(\comparator/N205 ) );
  xor2 \comparator/C1135  ( .a(a[919]), .b(b[919]), .out(\comparator/N207 ) );
  xor2 \comparator/C1136  ( .a(a[918]), .b(b[918]), .out(\comparator/N209 ) );
  xor2 \comparator/C1137  ( .a(a[917]), .b(b[917]), .out(\comparator/N211 ) );
  xor2 \comparator/C1138  ( .a(a[916]), .b(b[916]), .out(\comparator/N213 ) );
  xor2 \comparator/C1139  ( .a(a[915]), .b(b[915]), .out(\comparator/N215 ) );
  xor2 \comparator/C1140  ( .a(a[914]), .b(b[914]), .out(\comparator/N217 ) );
  xor2 \comparator/C1141  ( .a(a[913]), .b(b[913]), .out(\comparator/N219 ) );
  xor2 \comparator/C1142  ( .a(a[912]), .b(b[912]), .out(\comparator/N221 ) );
  xor2 \comparator/C1143  ( .a(a[911]), .b(b[911]), .out(\comparator/N223 ) );
  xor2 \comparator/C1144  ( .a(a[910]), .b(b[910]), .out(\comparator/N225 ) );
  xor2 \comparator/C1145  ( .a(a[909]), .b(b[909]), .out(\comparator/N227 ) );
  xor2 \comparator/C1146  ( .a(a[908]), .b(b[908]), .out(\comparator/N229 ) );
  xor2 \comparator/C1147  ( .a(a[907]), .b(b[907]), .out(\comparator/N231 ) );
  xor2 \comparator/C1148  ( .a(a[906]), .b(b[906]), .out(\comparator/N233 ) );
  xor2 \comparator/C1149  ( .a(a[905]), .b(b[905]), .out(\comparator/N235 ) );
  xor2 \comparator/C1150  ( .a(a[904]), .b(b[904]), .out(\comparator/N237 ) );
  xor2 \comparator/C1151  ( .a(a[903]), .b(b[903]), .out(\comparator/N239 ) );
  xor2 \comparator/C1152  ( .a(a[902]), .b(b[902]), .out(\comparator/N241 ) );
  xor2 \comparator/C1153  ( .a(a[901]), .b(b[901]), .out(\comparator/N243 ) );
  xor2 \comparator/C1154  ( .a(a[900]), .b(b[900]), .out(\comparator/N245 ) );
  xor2 \comparator/C1155  ( .a(a[899]), .b(b[899]), .out(\comparator/N247 ) );
  xor2 \comparator/C1156  ( .a(a[898]), .b(b[898]), .out(\comparator/N249 ) );
  xor2 \comparator/C1157  ( .a(a[897]), .b(b[897]), .out(\comparator/N251 ) );
  xor2 \comparator/C1158  ( .a(a[896]), .b(b[896]), .out(\comparator/N253 ) );
  xor2 \comparator/C1159  ( .a(a[895]), .b(b[895]), .out(\comparator/N255 ) );
  xor2 \comparator/C1160  ( .a(a[894]), .b(b[894]), .out(\comparator/N257 ) );
  xor2 \comparator/C1161  ( .a(a[893]), .b(b[893]), .out(\comparator/N259 ) );
  xor2 \comparator/C1162  ( .a(a[892]), .b(b[892]), .out(\comparator/N261 ) );
  xor2 \comparator/C1163  ( .a(a[891]), .b(b[891]), .out(\comparator/N263 ) );
  xor2 \comparator/C1164  ( .a(a[890]), .b(b[890]), .out(\comparator/N265 ) );
  xor2 \comparator/C1165  ( .a(a[889]), .b(b[889]), .out(\comparator/N267 ) );
  xor2 \comparator/C1166  ( .a(a[888]), .b(b[888]), .out(\comparator/N269 ) );
  xor2 \comparator/C1167  ( .a(a[887]), .b(b[887]), .out(\comparator/N271 ) );
  xor2 \comparator/C1168  ( .a(a[886]), .b(b[886]), .out(\comparator/N273 ) );
  xor2 \comparator/C1169  ( .a(a[885]), .b(b[885]), .out(\comparator/N275 ) );
  xor2 \comparator/C1170  ( .a(a[884]), .b(b[884]), .out(\comparator/N277 ) );
  xor2 \comparator/C1171  ( .a(a[883]), .b(b[883]), .out(\comparator/N279 ) );
  xor2 \comparator/C1172  ( .a(a[882]), .b(b[882]), .out(\comparator/N281 ) );
  xor2 \comparator/C1173  ( .a(a[881]), .b(b[881]), .out(\comparator/N283 ) );
  xor2 \comparator/C1174  ( .a(a[880]), .b(b[880]), .out(\comparator/N285 ) );
  xor2 \comparator/C1175  ( .a(a[879]), .b(b[879]), .out(\comparator/N287 ) );
  xor2 \comparator/C1176  ( .a(a[878]), .b(b[878]), .out(\comparator/N289 ) );
  xor2 \comparator/C1177  ( .a(a[877]), .b(b[877]), .out(\comparator/N291 ) );
  xor2 \comparator/C1178  ( .a(a[876]), .b(b[876]), .out(\comparator/N293 ) );
  xor2 \comparator/C1179  ( .a(a[875]), .b(b[875]), .out(\comparator/N295 ) );
  xor2 \comparator/C1180  ( .a(a[874]), .b(b[874]), .out(\comparator/N297 ) );
  xor2 \comparator/C1181  ( .a(a[873]), .b(b[873]), .out(\comparator/N299 ) );
  xor2 \comparator/C1182  ( .a(a[872]), .b(b[872]), .out(\comparator/N301 ) );
  xor2 \comparator/C1183  ( .a(a[871]), .b(b[871]), .out(\comparator/N303 ) );
  xor2 \comparator/C1184  ( .a(a[870]), .b(b[870]), .out(\comparator/N305 ) );
  xor2 \comparator/C1185  ( .a(a[869]), .b(b[869]), .out(\comparator/N307 ) );
  xor2 \comparator/C1186  ( .a(a[868]), .b(b[868]), .out(\comparator/N309 ) );
  xor2 \comparator/C1187  ( .a(a[867]), .b(b[867]), .out(\comparator/N311 ) );
  xor2 \comparator/C1188  ( .a(a[866]), .b(b[866]), .out(\comparator/N313 ) );
  xor2 \comparator/C1189  ( .a(a[865]), .b(b[865]), .out(\comparator/N315 ) );
  xor2 \comparator/C1190  ( .a(a[864]), .b(b[864]), .out(\comparator/N317 ) );
  xor2 \comparator/C1191  ( .a(a[863]), .b(b[863]), .out(\comparator/N319 ) );
  xor2 \comparator/C1192  ( .a(a[862]), .b(b[862]), .out(\comparator/N321 ) );
  xor2 \comparator/C1193  ( .a(a[861]), .b(b[861]), .out(\comparator/N323 ) );
  xor2 \comparator/C1194  ( .a(a[860]), .b(b[860]), .out(\comparator/N325 ) );
  xor2 \comparator/C1195  ( .a(a[859]), .b(b[859]), .out(\comparator/N327 ) );
  xor2 \comparator/C1196  ( .a(a[858]), .b(b[858]), .out(\comparator/N329 ) );
  xor2 \comparator/C1197  ( .a(a[857]), .b(b[857]), .out(\comparator/N331 ) );
  xor2 \comparator/C1198  ( .a(a[856]), .b(b[856]), .out(\comparator/N333 ) );
  xor2 \comparator/C1199  ( .a(a[855]), .b(b[855]), .out(\comparator/N335 ) );
  xor2 \comparator/C1200  ( .a(a[854]), .b(b[854]), .out(\comparator/N337 ) );
  xor2 \comparator/C1201  ( .a(a[853]), .b(b[853]), .out(\comparator/N339 ) );
  xor2 \comparator/C1202  ( .a(a[852]), .b(b[852]), .out(\comparator/N341 ) );
  xor2 \comparator/C1203  ( .a(a[851]), .b(b[851]), .out(\comparator/N343 ) );
  xor2 \comparator/C1204  ( .a(a[850]), .b(b[850]), .out(\comparator/N345 ) );
  xor2 \comparator/C1205  ( .a(a[849]), .b(b[849]), .out(\comparator/N347 ) );
  xor2 \comparator/C1206  ( .a(a[848]), .b(b[848]), .out(\comparator/N349 ) );
  xor2 \comparator/C1207  ( .a(a[847]), .b(b[847]), .out(\comparator/N351 ) );
  xor2 \comparator/C1208  ( .a(a[846]), .b(b[846]), .out(\comparator/N353 ) );
  xor2 \comparator/C1209  ( .a(a[845]), .b(b[845]), .out(\comparator/N355 ) );
  xor2 \comparator/C1210  ( .a(a[844]), .b(b[844]), .out(\comparator/N357 ) );
  xor2 \comparator/C1211  ( .a(a[843]), .b(b[843]), .out(\comparator/N359 ) );
  xor2 \comparator/C1212  ( .a(a[842]), .b(b[842]), .out(\comparator/N361 ) );
  xor2 \comparator/C1213  ( .a(a[841]), .b(b[841]), .out(\comparator/N363 ) );
  xor2 \comparator/C1214  ( .a(a[840]), .b(b[840]), .out(\comparator/N365 ) );
  xor2 \comparator/C1215  ( .a(a[839]), .b(b[839]), .out(\comparator/N367 ) );
  xor2 \comparator/C1216  ( .a(a[838]), .b(b[838]), .out(\comparator/N369 ) );
  xor2 \comparator/C1217  ( .a(a[837]), .b(b[837]), .out(\comparator/N371 ) );
  xor2 \comparator/C1218  ( .a(a[836]), .b(b[836]), .out(\comparator/N373 ) );
  xor2 \comparator/C1219  ( .a(a[835]), .b(b[835]), .out(\comparator/N375 ) );
  xor2 \comparator/C1220  ( .a(a[834]), .b(b[834]), .out(\comparator/N377 ) );
  xor2 \comparator/C1221  ( .a(a[833]), .b(b[833]), .out(\comparator/N379 ) );
  xor2 \comparator/C1222  ( .a(a[832]), .b(b[832]), .out(\comparator/N381 ) );
  xor2 \comparator/C1223  ( .a(a[831]), .b(b[831]), .out(\comparator/N383 ) );
  xor2 \comparator/C1224  ( .a(a[830]), .b(b[830]), .out(\comparator/N385 ) );
  xor2 \comparator/C1225  ( .a(a[829]), .b(b[829]), .out(\comparator/N387 ) );
  xor2 \comparator/C1226  ( .a(a[828]), .b(b[828]), .out(\comparator/N389 ) );
  xor2 \comparator/C1227  ( .a(a[827]), .b(b[827]), .out(\comparator/N391 ) );
  xor2 \comparator/C1228  ( .a(a[826]), .b(b[826]), .out(\comparator/N393 ) );
  xor2 \comparator/C1229  ( .a(a[825]), .b(b[825]), .out(\comparator/N395 ) );
  xor2 \comparator/C1230  ( .a(a[824]), .b(b[824]), .out(\comparator/N397 ) );
  xor2 \comparator/C1231  ( .a(a[823]), .b(b[823]), .out(\comparator/N399 ) );
  xor2 \comparator/C1232  ( .a(a[822]), .b(b[822]), .out(\comparator/N401 ) );
  xor2 \comparator/C1233  ( .a(a[821]), .b(b[821]), .out(\comparator/N403 ) );
  xor2 \comparator/C1234  ( .a(a[820]), .b(b[820]), .out(\comparator/N405 ) );
  xor2 \comparator/C1235  ( .a(a[819]), .b(b[819]), .out(\comparator/N407 ) );
  xor2 \comparator/C1236  ( .a(a[818]), .b(b[818]), .out(\comparator/N409 ) );
  xor2 \comparator/C1237  ( .a(a[817]), .b(b[817]), .out(\comparator/N411 ) );
  xor2 \comparator/C1238  ( .a(a[816]), .b(b[816]), .out(\comparator/N413 ) );
  xor2 \comparator/C1239  ( .a(a[815]), .b(b[815]), .out(\comparator/N415 ) );
  xor2 \comparator/C1240  ( .a(a[814]), .b(b[814]), .out(\comparator/N417 ) );
  xor2 \comparator/C1241  ( .a(a[813]), .b(b[813]), .out(\comparator/N419 ) );
  xor2 \comparator/C1242  ( .a(a[812]), .b(b[812]), .out(\comparator/N421 ) );
  xor2 \comparator/C1243  ( .a(a[811]), .b(b[811]), .out(\comparator/N423 ) );
  xor2 \comparator/C1244  ( .a(a[810]), .b(b[810]), .out(\comparator/N425 ) );
  xor2 \comparator/C1245  ( .a(a[809]), .b(b[809]), .out(\comparator/N427 ) );
  xor2 \comparator/C1246  ( .a(a[808]), .b(b[808]), .out(\comparator/N429 ) );
  xor2 \comparator/C1247  ( .a(a[807]), .b(b[807]), .out(\comparator/N431 ) );
  xor2 \comparator/C1248  ( .a(a[806]), .b(b[806]), .out(\comparator/N433 ) );
  xor2 \comparator/C1249  ( .a(a[805]), .b(b[805]), .out(\comparator/N435 ) );
  xor2 \comparator/C1250  ( .a(a[804]), .b(b[804]), .out(\comparator/N437 ) );
  xor2 \comparator/C1251  ( .a(a[803]), .b(b[803]), .out(\comparator/N439 ) );
  xor2 \comparator/C1252  ( .a(a[802]), .b(b[802]), .out(\comparator/N441 ) );
  xor2 \comparator/C1253  ( .a(a[801]), .b(b[801]), .out(\comparator/N443 ) );
  xor2 \comparator/C1254  ( .a(a[800]), .b(b[800]), .out(\comparator/N445 ) );
  xor2 \comparator/C1255  ( .a(a[799]), .b(b[799]), .out(\comparator/N447 ) );
  xor2 \comparator/C1256  ( .a(a[798]), .b(b[798]), .out(\comparator/N449 ) );
  xor2 \comparator/C1257  ( .a(a[797]), .b(b[797]), .out(\comparator/N451 ) );
  xor2 \comparator/C1258  ( .a(a[796]), .b(b[796]), .out(\comparator/N453 ) );
  xor2 \comparator/C1259  ( .a(a[795]), .b(b[795]), .out(\comparator/N455 ) );
  xor2 \comparator/C1260  ( .a(a[794]), .b(b[794]), .out(\comparator/N457 ) );
  xor2 \comparator/C1261  ( .a(a[793]), .b(b[793]), .out(\comparator/N459 ) );
  xor2 \comparator/C1262  ( .a(a[792]), .b(b[792]), .out(\comparator/N461 ) );
  xor2 \comparator/C1263  ( .a(a[791]), .b(b[791]), .out(\comparator/N463 ) );
  xor2 \comparator/C1264  ( .a(a[790]), .b(b[790]), .out(\comparator/N465 ) );
  xor2 \comparator/C1265  ( .a(a[789]), .b(b[789]), .out(\comparator/N467 ) );
  xor2 \comparator/C1266  ( .a(a[788]), .b(b[788]), .out(\comparator/N469 ) );
  xor2 \comparator/C1267  ( .a(a[787]), .b(b[787]), .out(\comparator/N471 ) );
  xor2 \comparator/C1268  ( .a(a[786]), .b(b[786]), .out(\comparator/N473 ) );
  xor2 \comparator/C1269  ( .a(a[785]), .b(b[785]), .out(\comparator/N475 ) );
  xor2 \comparator/C1270  ( .a(a[784]), .b(b[784]), .out(\comparator/N477 ) );
  xor2 \comparator/C1271  ( .a(a[783]), .b(b[783]), .out(\comparator/N479 ) );
  xor2 \comparator/C1272  ( .a(a[782]), .b(b[782]), .out(\comparator/N481 ) );
  xor2 \comparator/C1273  ( .a(a[781]), .b(b[781]), .out(\comparator/N483 ) );
  xor2 \comparator/C1274  ( .a(a[780]), .b(b[780]), .out(\comparator/N485 ) );
  xor2 \comparator/C1275  ( .a(a[779]), .b(b[779]), .out(\comparator/N487 ) );
  xor2 \comparator/C1276  ( .a(a[778]), .b(b[778]), .out(\comparator/N489 ) );
  xor2 \comparator/C1277  ( .a(a[777]), .b(b[777]), .out(\comparator/N491 ) );
  xor2 \comparator/C1278  ( .a(a[776]), .b(b[776]), .out(\comparator/N493 ) );
  xor2 \comparator/C1279  ( .a(a[775]), .b(b[775]), .out(\comparator/N495 ) );
  xor2 \comparator/C1280  ( .a(a[774]), .b(b[774]), .out(\comparator/N497 ) );
  xor2 \comparator/C1281  ( .a(a[773]), .b(b[773]), .out(\comparator/N499 ) );
  xor2 \comparator/C1282  ( .a(a[772]), .b(b[772]), .out(\comparator/N501 ) );
  xor2 \comparator/C1283  ( .a(a[771]), .b(b[771]), .out(\comparator/N503 ) );
  xor2 \comparator/C1284  ( .a(a[770]), .b(b[770]), .out(\comparator/N505 ) );
  xor2 \comparator/C1285  ( .a(a[769]), .b(b[769]), .out(\comparator/N507 ) );
  xor2 \comparator/C1286  ( .a(a[768]), .b(b[768]), .out(\comparator/N509 ) );
  xor2 \comparator/C1287  ( .a(a[767]), .b(b[767]), .out(\comparator/N511 ) );
  xor2 \comparator/C1288  ( .a(a[766]), .b(b[766]), .out(\comparator/N513 ) );
  xor2 \comparator/C1289  ( .a(a[765]), .b(b[765]), .out(\comparator/N515 ) );
  xor2 \comparator/C1290  ( .a(a[764]), .b(b[764]), .out(\comparator/N517 ) );
  xor2 \comparator/C1291  ( .a(a[763]), .b(b[763]), .out(\comparator/N519 ) );
  xor2 \comparator/C1292  ( .a(a[762]), .b(b[762]), .out(\comparator/N521 ) );
  xor2 \comparator/C1293  ( .a(a[761]), .b(b[761]), .out(\comparator/N523 ) );
  xor2 \comparator/C1294  ( .a(a[760]), .b(b[760]), .out(\comparator/N525 ) );
  xor2 \comparator/C1295  ( .a(a[759]), .b(b[759]), .out(\comparator/N527 ) );
  xor2 \comparator/C1296  ( .a(a[758]), .b(b[758]), .out(\comparator/N529 ) );
  xor2 \comparator/C1297  ( .a(a[757]), .b(b[757]), .out(\comparator/N531 ) );
  xor2 \comparator/C1298  ( .a(a[756]), .b(b[756]), .out(\comparator/N533 ) );
  xor2 \comparator/C1299  ( .a(a[755]), .b(b[755]), .out(\comparator/N535 ) );
  xor2 \comparator/C1300  ( .a(a[754]), .b(b[754]), .out(\comparator/N537 ) );
  xor2 \comparator/C1301  ( .a(a[753]), .b(b[753]), .out(\comparator/N539 ) );
  xor2 \comparator/C1302  ( .a(a[752]), .b(b[752]), .out(\comparator/N541 ) );
  xor2 \comparator/C1303  ( .a(a[751]), .b(b[751]), .out(\comparator/N543 ) );
  xor2 \comparator/C1304  ( .a(a[750]), .b(b[750]), .out(\comparator/N545 ) );
  xor2 \comparator/C1305  ( .a(a[749]), .b(b[749]), .out(\comparator/N547 ) );
  xor2 \comparator/C1306  ( .a(a[748]), .b(b[748]), .out(\comparator/N549 ) );
  xor2 \comparator/C1307  ( .a(a[747]), .b(b[747]), .out(\comparator/N551 ) );
  xor2 \comparator/C1308  ( .a(a[746]), .b(b[746]), .out(\comparator/N553 ) );
  xor2 \comparator/C1309  ( .a(a[745]), .b(b[745]), .out(\comparator/N555 ) );
  xor2 \comparator/C1310  ( .a(a[744]), .b(b[744]), .out(\comparator/N557 ) );
  xor2 \comparator/C1311  ( .a(a[743]), .b(b[743]), .out(\comparator/N559 ) );
  xor2 \comparator/C1312  ( .a(a[742]), .b(b[742]), .out(\comparator/N561 ) );
  xor2 \comparator/C1313  ( .a(a[741]), .b(b[741]), .out(\comparator/N563 ) );
  xor2 \comparator/C1314  ( .a(a[740]), .b(b[740]), .out(\comparator/N565 ) );
  xor2 \comparator/C1315  ( .a(a[739]), .b(b[739]), .out(\comparator/N567 ) );
  xor2 \comparator/C1316  ( .a(a[738]), .b(b[738]), .out(\comparator/N569 ) );
  xor2 \comparator/C1317  ( .a(a[737]), .b(b[737]), .out(\comparator/N571 ) );
  xor2 \comparator/C1318  ( .a(a[736]), .b(b[736]), .out(\comparator/N573 ) );
  xor2 \comparator/C1319  ( .a(a[735]), .b(b[735]), .out(\comparator/N575 ) );
  xor2 \comparator/C1320  ( .a(a[734]), .b(b[734]), .out(\comparator/N577 ) );
  xor2 \comparator/C1321  ( .a(a[733]), .b(b[733]), .out(\comparator/N579 ) );
  xor2 \comparator/C1322  ( .a(a[732]), .b(b[732]), .out(\comparator/N581 ) );
  xor2 \comparator/C1323  ( .a(a[731]), .b(b[731]), .out(\comparator/N583 ) );
  xor2 \comparator/C1324  ( .a(a[730]), .b(b[730]), .out(\comparator/N585 ) );
  xor2 \comparator/C1325  ( .a(a[729]), .b(b[729]), .out(\comparator/N587 ) );
  xor2 \comparator/C1326  ( .a(a[728]), .b(b[728]), .out(\comparator/N589 ) );
  xor2 \comparator/C1327  ( .a(a[727]), .b(b[727]), .out(\comparator/N591 ) );
  xor2 \comparator/C1328  ( .a(a[726]), .b(b[726]), .out(\comparator/N593 ) );
  xor2 \comparator/C1329  ( .a(a[725]), .b(b[725]), .out(\comparator/N595 ) );
  xor2 \comparator/C1330  ( .a(a[724]), .b(b[724]), .out(\comparator/N597 ) );
  xor2 \comparator/C1331  ( .a(a[723]), .b(b[723]), .out(\comparator/N599 ) );
  xor2 \comparator/C1332  ( .a(a[722]), .b(b[722]), .out(\comparator/N601 ) );
  xor2 \comparator/C1333  ( .a(a[721]), .b(b[721]), .out(\comparator/N603 ) );
  xor2 \comparator/C1334  ( .a(a[720]), .b(b[720]), .out(\comparator/N605 ) );
  xor2 \comparator/C1335  ( .a(a[719]), .b(b[719]), .out(\comparator/N607 ) );
  xor2 \comparator/C1336  ( .a(a[718]), .b(b[718]), .out(\comparator/N609 ) );
  xor2 \comparator/C1337  ( .a(a[717]), .b(b[717]), .out(\comparator/N611 ) );
  xor2 \comparator/C1338  ( .a(a[716]), .b(b[716]), .out(\comparator/N613 ) );
  xor2 \comparator/C1339  ( .a(a[715]), .b(b[715]), .out(\comparator/N615 ) );
  xor2 \comparator/C1340  ( .a(a[714]), .b(b[714]), .out(\comparator/N617 ) );
  xor2 \comparator/C1341  ( .a(a[713]), .b(b[713]), .out(\comparator/N619 ) );
  xor2 \comparator/C1342  ( .a(a[712]), .b(b[712]), .out(\comparator/N621 ) );
  xor2 \comparator/C1343  ( .a(a[711]), .b(b[711]), .out(\comparator/N623 ) );
  xor2 \comparator/C1344  ( .a(a[710]), .b(b[710]), .out(\comparator/N625 ) );
  xor2 \comparator/C1345  ( .a(a[709]), .b(b[709]), .out(\comparator/N627 ) );
  xor2 \comparator/C1346  ( .a(a[708]), .b(b[708]), .out(\comparator/N629 ) );
  xor2 \comparator/C1347  ( .a(a[707]), .b(b[707]), .out(\comparator/N631 ) );
  xor2 \comparator/C1348  ( .a(a[706]), .b(b[706]), .out(\comparator/N633 ) );
  xor2 \comparator/C1349  ( .a(a[705]), .b(b[705]), .out(\comparator/N635 ) );
  xor2 \comparator/C1350  ( .a(a[704]), .b(b[704]), .out(\comparator/N637 ) );
  xor2 \comparator/C1351  ( .a(a[703]), .b(b[703]), .out(\comparator/N639 ) );
  xor2 \comparator/C1352  ( .a(a[702]), .b(b[702]), .out(\comparator/N641 ) );
  xor2 \comparator/C1353  ( .a(a[701]), .b(b[701]), .out(\comparator/N643 ) );
  xor2 \comparator/C1354  ( .a(a[700]), .b(b[700]), .out(\comparator/N645 ) );
  xor2 \comparator/C1355  ( .a(a[699]), .b(b[699]), .out(\comparator/N647 ) );
  xor2 \comparator/C1356  ( .a(a[698]), .b(b[698]), .out(\comparator/N649 ) );
  xor2 \comparator/C1357  ( .a(a[697]), .b(b[697]), .out(\comparator/N651 ) );
  xor2 \comparator/C1358  ( .a(a[696]), .b(b[696]), .out(\comparator/N653 ) );
  xor2 \comparator/C1359  ( .a(a[695]), .b(b[695]), .out(\comparator/N655 ) );
  xor2 \comparator/C1360  ( .a(a[694]), .b(b[694]), .out(\comparator/N657 ) );
  xor2 \comparator/C1361  ( .a(a[693]), .b(b[693]), .out(\comparator/N659 ) );
  xor2 \comparator/C1362  ( .a(a[692]), .b(b[692]), .out(\comparator/N661 ) );
  xor2 \comparator/C1363  ( .a(a[691]), .b(b[691]), .out(\comparator/N663 ) );
  xor2 \comparator/C1364  ( .a(a[690]), .b(b[690]), .out(\comparator/N665 ) );
  xor2 \comparator/C1365  ( .a(a[689]), .b(b[689]), .out(\comparator/N667 ) );
  xor2 \comparator/C1366  ( .a(a[688]), .b(b[688]), .out(\comparator/N669 ) );
  xor2 \comparator/C1367  ( .a(a[687]), .b(b[687]), .out(\comparator/N671 ) );
  xor2 \comparator/C1368  ( .a(a[686]), .b(b[686]), .out(\comparator/N673 ) );
  xor2 \comparator/C1369  ( .a(a[685]), .b(b[685]), .out(\comparator/N675 ) );
  xor2 \comparator/C1370  ( .a(a[684]), .b(b[684]), .out(\comparator/N677 ) );
  xor2 \comparator/C1371  ( .a(a[683]), .b(b[683]), .out(\comparator/N679 ) );
  xor2 \comparator/C1372  ( .a(a[682]), .b(b[682]), .out(\comparator/N681 ) );
  xor2 \comparator/C1373  ( .a(a[681]), .b(b[681]), .out(\comparator/N683 ) );
  xor2 \comparator/C1374  ( .a(a[680]), .b(b[680]), .out(\comparator/N685 ) );
  xor2 \comparator/C1375  ( .a(a[679]), .b(b[679]), .out(\comparator/N687 ) );
  xor2 \comparator/C1376  ( .a(a[678]), .b(b[678]), .out(\comparator/N689 ) );
  xor2 \comparator/C1377  ( .a(a[677]), .b(b[677]), .out(\comparator/N691 ) );
  xor2 \comparator/C1378  ( .a(a[676]), .b(b[676]), .out(\comparator/N693 ) );
  xor2 \comparator/C1379  ( .a(a[675]), .b(b[675]), .out(\comparator/N695 ) );
  xor2 \comparator/C1380  ( .a(a[674]), .b(b[674]), .out(\comparator/N697 ) );
  xor2 \comparator/C1381  ( .a(a[673]), .b(b[673]), .out(\comparator/N699 ) );
  xor2 \comparator/C1382  ( .a(a[672]), .b(b[672]), .out(\comparator/N701 ) );
  xor2 \comparator/C1383  ( .a(a[671]), .b(b[671]), .out(\comparator/N703 ) );
  xor2 \comparator/C1384  ( .a(a[670]), .b(b[670]), .out(\comparator/N705 ) );
  xor2 \comparator/C1385  ( .a(a[669]), .b(b[669]), .out(\comparator/N707 ) );
  xor2 \comparator/C1386  ( .a(a[668]), .b(b[668]), .out(\comparator/N709 ) );
  xor2 \comparator/C1387  ( .a(a[667]), .b(b[667]), .out(\comparator/N711 ) );
  xor2 \comparator/C1388  ( .a(a[666]), .b(b[666]), .out(\comparator/N713 ) );
  xor2 \comparator/C1389  ( .a(a[665]), .b(b[665]), .out(\comparator/N715 ) );
  xor2 \comparator/C1390  ( .a(a[664]), .b(b[664]), .out(\comparator/N717 ) );
  xor2 \comparator/C1391  ( .a(a[663]), .b(b[663]), .out(\comparator/N719 ) );
  xor2 \comparator/C1392  ( .a(a[662]), .b(b[662]), .out(\comparator/N721 ) );
  xor2 \comparator/C1393  ( .a(a[661]), .b(b[661]), .out(\comparator/N723 ) );
  xor2 \comparator/C1394  ( .a(a[660]), .b(b[660]), .out(\comparator/N725 ) );
  xor2 \comparator/C1395  ( .a(a[659]), .b(b[659]), .out(\comparator/N727 ) );
  xor2 \comparator/C1396  ( .a(a[658]), .b(b[658]), .out(\comparator/N729 ) );
  xor2 \comparator/C1397  ( .a(a[657]), .b(b[657]), .out(\comparator/N731 ) );
  xor2 \comparator/C1398  ( .a(a[656]), .b(b[656]), .out(\comparator/N733 ) );
  xor2 \comparator/C1399  ( .a(a[655]), .b(b[655]), .out(\comparator/N735 ) );
  xor2 \comparator/C1400  ( .a(a[654]), .b(b[654]), .out(\comparator/N737 ) );
  xor2 \comparator/C1401  ( .a(a[653]), .b(b[653]), .out(\comparator/N739 ) );
  xor2 \comparator/C1402  ( .a(a[652]), .b(b[652]), .out(\comparator/N741 ) );
  xor2 \comparator/C1403  ( .a(a[651]), .b(b[651]), .out(\comparator/N743 ) );
  xor2 \comparator/C1404  ( .a(a[650]), .b(b[650]), .out(\comparator/N745 ) );
  xor2 \comparator/C1405  ( .a(a[649]), .b(b[649]), .out(\comparator/N747 ) );
  xor2 \comparator/C1406  ( .a(a[648]), .b(b[648]), .out(\comparator/N749 ) );
  xor2 \comparator/C1407  ( .a(a[647]), .b(b[647]), .out(\comparator/N751 ) );
  xor2 \comparator/C1408  ( .a(a[646]), .b(b[646]), .out(\comparator/N753 ) );
  xor2 \comparator/C1409  ( .a(a[645]), .b(b[645]), .out(\comparator/N755 ) );
  xor2 \comparator/C1410  ( .a(a[644]), .b(b[644]), .out(\comparator/N757 ) );
  xor2 \comparator/C1411  ( .a(a[643]), .b(b[643]), .out(\comparator/N759 ) );
  xor2 \comparator/C1412  ( .a(a[642]), .b(b[642]), .out(\comparator/N761 ) );
  xor2 \comparator/C1413  ( .a(a[641]), .b(b[641]), .out(\comparator/N763 ) );
  xor2 \comparator/C1414  ( .a(a[640]), .b(b[640]), .out(\comparator/N765 ) );
  xor2 \comparator/C1415  ( .a(a[639]), .b(b[639]), .out(\comparator/N767 ) );
  xor2 \comparator/C1416  ( .a(a[638]), .b(b[638]), .out(\comparator/N769 ) );
  xor2 \comparator/C1417  ( .a(a[637]), .b(b[637]), .out(\comparator/N771 ) );
  xor2 \comparator/C1418  ( .a(a[636]), .b(b[636]), .out(\comparator/N773 ) );
  xor2 \comparator/C1419  ( .a(a[635]), .b(b[635]), .out(\comparator/N775 ) );
  xor2 \comparator/C1420  ( .a(a[634]), .b(b[634]), .out(\comparator/N777 ) );
  xor2 \comparator/C1421  ( .a(a[633]), .b(b[633]), .out(\comparator/N779 ) );
  xor2 \comparator/C1422  ( .a(a[632]), .b(b[632]), .out(\comparator/N781 ) );
  xor2 \comparator/C1423  ( .a(a[631]), .b(b[631]), .out(\comparator/N783 ) );
  xor2 \comparator/C1424  ( .a(a[630]), .b(b[630]), .out(\comparator/N785 ) );
  xor2 \comparator/C1425  ( .a(a[629]), .b(b[629]), .out(\comparator/N787 ) );
  xor2 \comparator/C1426  ( .a(a[628]), .b(b[628]), .out(\comparator/N789 ) );
  xor2 \comparator/C1427  ( .a(a[627]), .b(b[627]), .out(\comparator/N791 ) );
  xor2 \comparator/C1428  ( .a(a[626]), .b(b[626]), .out(\comparator/N793 ) );
  xor2 \comparator/C1429  ( .a(a[625]), .b(b[625]), .out(\comparator/N795 ) );
  xor2 \comparator/C1430  ( .a(a[624]), .b(b[624]), .out(\comparator/N797 ) );
  xor2 \comparator/C1431  ( .a(a[623]), .b(b[623]), .out(\comparator/N799 ) );
  xor2 \comparator/C1432  ( .a(a[622]), .b(b[622]), .out(\comparator/N801 ) );
  xor2 \comparator/C1433  ( .a(a[621]), .b(b[621]), .out(\comparator/N803 ) );
  xor2 \comparator/C1434  ( .a(a[620]), .b(b[620]), .out(\comparator/N805 ) );
  xor2 \comparator/C1435  ( .a(a[619]), .b(b[619]), .out(\comparator/N807 ) );
  xor2 \comparator/C1436  ( .a(a[618]), .b(b[618]), .out(\comparator/N809 ) );
  xor2 \comparator/C1437  ( .a(a[617]), .b(b[617]), .out(\comparator/N811 ) );
  xor2 \comparator/C1438  ( .a(a[616]), .b(b[616]), .out(\comparator/N813 ) );
  xor2 \comparator/C1439  ( .a(a[615]), .b(b[615]), .out(\comparator/N815 ) );
  xor2 \comparator/C1440  ( .a(a[614]), .b(b[614]), .out(\comparator/N817 ) );
  xor2 \comparator/C1441  ( .a(a[613]), .b(b[613]), .out(\comparator/N819 ) );
  xor2 \comparator/C1442  ( .a(a[612]), .b(b[612]), .out(\comparator/N821 ) );
  xor2 \comparator/C1443  ( .a(a[611]), .b(b[611]), .out(\comparator/N823 ) );
  xor2 \comparator/C1444  ( .a(a[610]), .b(b[610]), .out(\comparator/N825 ) );
  xor2 \comparator/C1445  ( .a(a[609]), .b(b[609]), .out(\comparator/N827 ) );
  xor2 \comparator/C1446  ( .a(a[608]), .b(b[608]), .out(\comparator/N829 ) );
  xor2 \comparator/C1447  ( .a(a[607]), .b(b[607]), .out(\comparator/N831 ) );
  xor2 \comparator/C1448  ( .a(a[606]), .b(b[606]), .out(\comparator/N833 ) );
  xor2 \comparator/C1449  ( .a(a[605]), .b(b[605]), .out(\comparator/N835 ) );
  xor2 \comparator/C1450  ( .a(a[604]), .b(b[604]), .out(\comparator/N837 ) );
  xor2 \comparator/C1451  ( .a(a[603]), .b(b[603]), .out(\comparator/N839 ) );
  xor2 \comparator/C1452  ( .a(a[602]), .b(b[602]), .out(\comparator/N841 ) );
  xor2 \comparator/C1453  ( .a(a[601]), .b(b[601]), .out(\comparator/N843 ) );
  xor2 \comparator/C1454  ( .a(a[600]), .b(b[600]), .out(\comparator/N845 ) );
  xor2 \comparator/C1455  ( .a(a[599]), .b(b[599]), .out(\comparator/N847 ) );
  xor2 \comparator/C1456  ( .a(a[598]), .b(b[598]), .out(\comparator/N849 ) );
  xor2 \comparator/C1457  ( .a(a[597]), .b(b[597]), .out(\comparator/N851 ) );
  xor2 \comparator/C1458  ( .a(a[596]), .b(b[596]), .out(\comparator/N853 ) );
  xor2 \comparator/C1459  ( .a(a[595]), .b(b[595]), .out(\comparator/N855 ) );
  xor2 \comparator/C1460  ( .a(a[594]), .b(b[594]), .out(\comparator/N857 ) );
  xor2 \comparator/C1461  ( .a(a[593]), .b(b[593]), .out(\comparator/N859 ) );
  xor2 \comparator/C1462  ( .a(a[592]), .b(b[592]), .out(\comparator/N861 ) );
  xor2 \comparator/C1463  ( .a(a[591]), .b(b[591]), .out(\comparator/N863 ) );
  xor2 \comparator/C1464  ( .a(a[590]), .b(b[590]), .out(\comparator/N865 ) );
  xor2 \comparator/C1465  ( .a(a[589]), .b(b[589]), .out(\comparator/N867 ) );
  xor2 \comparator/C1466  ( .a(a[588]), .b(b[588]), .out(\comparator/N869 ) );
  xor2 \comparator/C1467  ( .a(a[587]), .b(b[587]), .out(\comparator/N871 ) );
  xor2 \comparator/C1468  ( .a(a[586]), .b(b[586]), .out(\comparator/N873 ) );
  xor2 \comparator/C1469  ( .a(a[585]), .b(b[585]), .out(\comparator/N875 ) );
  xor2 \comparator/C1470  ( .a(a[584]), .b(b[584]), .out(\comparator/N877 ) );
  xor2 \comparator/C1471  ( .a(a[583]), .b(b[583]), .out(\comparator/N879 ) );
  xor2 \comparator/C1472  ( .a(a[582]), .b(b[582]), .out(\comparator/N881 ) );
  xor2 \comparator/C1473  ( .a(a[581]), .b(b[581]), .out(\comparator/N883 ) );
  xor2 \comparator/C1474  ( .a(a[580]), .b(b[580]), .out(\comparator/N885 ) );
  xor2 \comparator/C1475  ( .a(a[579]), .b(b[579]), .out(\comparator/N887 ) );
  xor2 \comparator/C1476  ( .a(a[578]), .b(b[578]), .out(\comparator/N889 ) );
  xor2 \comparator/C1477  ( .a(a[577]), .b(b[577]), .out(\comparator/N891 ) );
  xor2 \comparator/C1478  ( .a(a[576]), .b(b[576]), .out(\comparator/N893 ) );
  xor2 \comparator/C1479  ( .a(a[575]), .b(b[575]), .out(\comparator/N895 ) );
  xor2 \comparator/C1480  ( .a(a[574]), .b(b[574]), .out(\comparator/N897 ) );
  xor2 \comparator/C1481  ( .a(a[573]), .b(b[573]), .out(\comparator/N899 ) );
  xor2 \comparator/C1482  ( .a(a[572]), .b(b[572]), .out(\comparator/N901 ) );
  xor2 \comparator/C1483  ( .a(a[571]), .b(b[571]), .out(\comparator/N903 ) );
  xor2 \comparator/C1484  ( .a(a[570]), .b(b[570]), .out(\comparator/N905 ) );
  xor2 \comparator/C1485  ( .a(a[569]), .b(b[569]), .out(\comparator/N907 ) );
  xor2 \comparator/C1486  ( .a(a[568]), .b(b[568]), .out(\comparator/N909 ) );
  xor2 \comparator/C1487  ( .a(a[567]), .b(b[567]), .out(\comparator/N911 ) );
  xor2 \comparator/C1488  ( .a(a[566]), .b(b[566]), .out(\comparator/N913 ) );
  xor2 \comparator/C1489  ( .a(a[565]), .b(b[565]), .out(\comparator/N915 ) );
  xor2 \comparator/C1490  ( .a(a[564]), .b(b[564]), .out(\comparator/N917 ) );
  xor2 \comparator/C1491  ( .a(a[563]), .b(b[563]), .out(\comparator/N919 ) );
  xor2 \comparator/C1492  ( .a(a[562]), .b(b[562]), .out(\comparator/N921 ) );
  xor2 \comparator/C1493  ( .a(a[561]), .b(b[561]), .out(\comparator/N923 ) );
  xor2 \comparator/C1494  ( .a(a[560]), .b(b[560]), .out(\comparator/N925 ) );
  xor2 \comparator/C1495  ( .a(a[559]), .b(b[559]), .out(\comparator/N927 ) );
  xor2 \comparator/C1496  ( .a(a[558]), .b(b[558]), .out(\comparator/N929 ) );
  xor2 \comparator/C1497  ( .a(a[557]), .b(b[557]), .out(\comparator/N931 ) );
  xor2 \comparator/C1498  ( .a(a[556]), .b(b[556]), .out(\comparator/N933 ) );
  xor2 \comparator/C1499  ( .a(a[555]), .b(b[555]), .out(\comparator/N935 ) );
  xor2 \comparator/C1500  ( .a(a[554]), .b(b[554]), .out(\comparator/N937 ) );
  xor2 \comparator/C1501  ( .a(a[553]), .b(b[553]), .out(\comparator/N939 ) );
  xor2 \comparator/C1502  ( .a(a[552]), .b(b[552]), .out(\comparator/N941 ) );
  xor2 \comparator/C1503  ( .a(a[551]), .b(b[551]), .out(\comparator/N943 ) );
  xor2 \comparator/C1504  ( .a(a[550]), .b(b[550]), .out(\comparator/N945 ) );
  xor2 \comparator/C1505  ( .a(a[549]), .b(b[549]), .out(\comparator/N947 ) );
  xor2 \comparator/C1506  ( .a(a[548]), .b(b[548]), .out(\comparator/N949 ) );
  xor2 \comparator/C1507  ( .a(a[547]), .b(b[547]), .out(\comparator/N951 ) );
  xor2 \comparator/C1508  ( .a(a[546]), .b(b[546]), .out(\comparator/N953 ) );
  xor2 \comparator/C1509  ( .a(a[545]), .b(b[545]), .out(\comparator/N955 ) );
  xor2 \comparator/C1510  ( .a(a[544]), .b(b[544]), .out(\comparator/N957 ) );
  xor2 \comparator/C1511  ( .a(a[543]), .b(b[543]), .out(\comparator/N959 ) );
  xor2 \comparator/C1512  ( .a(a[542]), .b(b[542]), .out(\comparator/N961 ) );
  xor2 \comparator/C1513  ( .a(a[541]), .b(b[541]), .out(\comparator/N963 ) );
  xor2 \comparator/C1514  ( .a(a[540]), .b(b[540]), .out(\comparator/N965 ) );
  xor2 \comparator/C1515  ( .a(a[539]), .b(b[539]), .out(\comparator/N967 ) );
  xor2 \comparator/C1516  ( .a(a[538]), .b(b[538]), .out(\comparator/N969 ) );
  xor2 \comparator/C1517  ( .a(a[537]), .b(b[537]), .out(\comparator/N971 ) );
  xor2 \comparator/C1518  ( .a(a[536]), .b(b[536]), .out(\comparator/N973 ) );
  xor2 \comparator/C1519  ( .a(a[535]), .b(b[535]), .out(\comparator/N975 ) );
  xor2 \comparator/C1520  ( .a(a[534]), .b(b[534]), .out(\comparator/N977 ) );
  xor2 \comparator/C1521  ( .a(a[533]), .b(b[533]), .out(\comparator/N979 ) );
  xor2 \comparator/C1522  ( .a(a[532]), .b(b[532]), .out(\comparator/N981 ) );
  xor2 \comparator/C1523  ( .a(a[531]), .b(b[531]), .out(\comparator/N983 ) );
  xor2 \comparator/C1524  ( .a(a[530]), .b(b[530]), .out(\comparator/N985 ) );
  xor2 \comparator/C1525  ( .a(a[529]), .b(b[529]), .out(\comparator/N987 ) );
  xor2 \comparator/C1526  ( .a(a[528]), .b(b[528]), .out(\comparator/N989 ) );
  xor2 \comparator/C1527  ( .a(a[527]), .b(b[527]), .out(\comparator/N991 ) );
  xor2 \comparator/C1528  ( .a(a[526]), .b(b[526]), .out(\comparator/N993 ) );
  xor2 \comparator/C1529  ( .a(a[525]), .b(b[525]), .out(\comparator/N995 ) );
  xor2 \comparator/C1530  ( .a(a[524]), .b(b[524]), .out(\comparator/N997 ) );
  xor2 \comparator/C1531  ( .a(a[523]), .b(b[523]), .out(\comparator/N999 ) );
  xor2 \comparator/C1532  ( .a(a[522]), .b(b[522]), .out(\comparator/N1001 )
         );
  xor2 \comparator/C1533  ( .a(a[521]), .b(b[521]), .out(\comparator/N1003 )
         );
  xor2 \comparator/C1534  ( .a(a[520]), .b(b[520]), .out(\comparator/N1005 )
         );
  xor2 \comparator/C1535  ( .a(a[519]), .b(b[519]), .out(\comparator/N1007 )
         );
  xor2 \comparator/C1536  ( .a(a[518]), .b(b[518]), .out(\comparator/N1009 )
         );
  xor2 \comparator/C1537  ( .a(a[517]), .b(b[517]), .out(\comparator/N1011 )
         );
  xor2 \comparator/C1538  ( .a(a[516]), .b(b[516]), .out(\comparator/N1013 )
         );
  xor2 \comparator/C1539  ( .a(a[515]), .b(b[515]), .out(\comparator/N1015 )
         );
  xor2 \comparator/C1540  ( .a(a[514]), .b(b[514]), .out(\comparator/N1017 )
         );
  xor2 \comparator/C1541  ( .a(a[513]), .b(b[513]), .out(\comparator/N1019 )
         );
  xor2 \comparator/C1542  ( .a(a[512]), .b(b[512]), .out(\comparator/N1021 )
         );
  xor2 \comparator/C1543  ( .a(a[511]), .b(b[511]), .out(\comparator/N1023 )
         );
  xor2 \comparator/C1544  ( .a(a[510]), .b(b[510]), .out(\comparator/N1025 )
         );
  xor2 \comparator/C1545  ( .a(a[509]), .b(b[509]), .out(\comparator/N1027 )
         );
  xor2 \comparator/C1546  ( .a(a[508]), .b(b[508]), .out(\comparator/N1029 )
         );
  xor2 \comparator/C1547  ( .a(a[507]), .b(b[507]), .out(\comparator/N1031 )
         );
  xor2 \comparator/C1548  ( .a(a[506]), .b(b[506]), .out(\comparator/N1033 )
         );
  xor2 \comparator/C1549  ( .a(a[505]), .b(b[505]), .out(\comparator/N1035 )
         );
  xor2 \comparator/C1550  ( .a(a[504]), .b(b[504]), .out(\comparator/N1037 )
         );
  xor2 \comparator/C1551  ( .a(a[503]), .b(b[503]), .out(\comparator/N1039 )
         );
  xor2 \comparator/C1552  ( .a(a[502]), .b(b[502]), .out(\comparator/N1041 )
         );
  xor2 \comparator/C1553  ( .a(a[501]), .b(b[501]), .out(\comparator/N1043 )
         );
  xor2 \comparator/C1554  ( .a(a[500]), .b(b[500]), .out(\comparator/N1045 )
         );
  xor2 \comparator/C1555  ( .a(a[499]), .b(b[499]), .out(\comparator/N1047 )
         );
  xor2 \comparator/C1556  ( .a(a[498]), .b(b[498]), .out(\comparator/N1049 )
         );
  xor2 \comparator/C1557  ( .a(a[497]), .b(b[497]), .out(\comparator/N1051 )
         );
  xor2 \comparator/C1558  ( .a(a[496]), .b(b[496]), .out(\comparator/N1053 )
         );
  xor2 \comparator/C1559  ( .a(a[495]), .b(b[495]), .out(\comparator/N1055 )
         );
  xor2 \comparator/C1560  ( .a(a[494]), .b(b[494]), .out(\comparator/N1057 )
         );
  xor2 \comparator/C1561  ( .a(a[493]), .b(b[493]), .out(\comparator/N1059 )
         );
  xor2 \comparator/C1562  ( .a(a[492]), .b(b[492]), .out(\comparator/N1061 )
         );
  xor2 \comparator/C1563  ( .a(a[491]), .b(b[491]), .out(\comparator/N1063 )
         );
  xor2 \comparator/C1564  ( .a(a[490]), .b(b[490]), .out(\comparator/N1065 )
         );
  xor2 \comparator/C1565  ( .a(a[489]), .b(b[489]), .out(\comparator/N1067 )
         );
  xor2 \comparator/C1566  ( .a(a[488]), .b(b[488]), .out(\comparator/N1069 )
         );
  xor2 \comparator/C1567  ( .a(a[487]), .b(b[487]), .out(\comparator/N1071 )
         );
  xor2 \comparator/C1568  ( .a(a[486]), .b(b[486]), .out(\comparator/N1073 )
         );
  xor2 \comparator/C1569  ( .a(a[485]), .b(b[485]), .out(\comparator/N1075 )
         );
  xor2 \comparator/C1570  ( .a(a[484]), .b(b[484]), .out(\comparator/N1077 )
         );
  xor2 \comparator/C1571  ( .a(a[483]), .b(b[483]), .out(\comparator/N1079 )
         );
  xor2 \comparator/C1572  ( .a(a[482]), .b(b[482]), .out(\comparator/N1081 )
         );
  xor2 \comparator/C1573  ( .a(a[481]), .b(b[481]), .out(\comparator/N1083 )
         );
  xor2 \comparator/C1574  ( .a(a[480]), .b(b[480]), .out(\comparator/N1085 )
         );
  xor2 \comparator/C1575  ( .a(a[479]), .b(b[479]), .out(\comparator/N1087 )
         );
  xor2 \comparator/C1576  ( .a(a[478]), .b(b[478]), .out(\comparator/N1089 )
         );
  xor2 \comparator/C1577  ( .a(a[477]), .b(b[477]), .out(\comparator/N1091 )
         );
  xor2 \comparator/C1578  ( .a(a[476]), .b(b[476]), .out(\comparator/N1093 )
         );
  xor2 \comparator/C1579  ( .a(a[475]), .b(b[475]), .out(\comparator/N1095 )
         );
  xor2 \comparator/C1580  ( .a(a[474]), .b(b[474]), .out(\comparator/N1097 )
         );
  xor2 \comparator/C1581  ( .a(a[473]), .b(b[473]), .out(\comparator/N1099 )
         );
  xor2 \comparator/C1582  ( .a(a[472]), .b(b[472]), .out(\comparator/N1101 )
         );
  xor2 \comparator/C1583  ( .a(a[471]), .b(b[471]), .out(\comparator/N1103 )
         );
  xor2 \comparator/C1584  ( .a(a[470]), .b(b[470]), .out(\comparator/N1105 )
         );
  xor2 \comparator/C1585  ( .a(a[469]), .b(b[469]), .out(\comparator/N1107 )
         );
  xor2 \comparator/C1586  ( .a(a[468]), .b(b[468]), .out(\comparator/N1109 )
         );
  xor2 \comparator/C1587  ( .a(a[467]), .b(b[467]), .out(\comparator/N1111 )
         );
  xor2 \comparator/C1588  ( .a(a[466]), .b(b[466]), .out(\comparator/N1113 )
         );
  xor2 \comparator/C1589  ( .a(a[465]), .b(b[465]), .out(\comparator/N1115 )
         );
  xor2 \comparator/C1590  ( .a(a[464]), .b(b[464]), .out(\comparator/N1117 )
         );
  xor2 \comparator/C1591  ( .a(a[463]), .b(b[463]), .out(\comparator/N1119 )
         );
  xor2 \comparator/C1592  ( .a(a[462]), .b(b[462]), .out(\comparator/N1121 )
         );
  xor2 \comparator/C1593  ( .a(a[461]), .b(b[461]), .out(\comparator/N1123 )
         );
  xor2 \comparator/C1594  ( .a(a[460]), .b(b[460]), .out(\comparator/N1125 )
         );
  xor2 \comparator/C1595  ( .a(a[459]), .b(b[459]), .out(\comparator/N1127 )
         );
  xor2 \comparator/C1596  ( .a(a[458]), .b(b[458]), .out(\comparator/N1129 )
         );
  xor2 \comparator/C1597  ( .a(a[457]), .b(b[457]), .out(\comparator/N1131 )
         );
  xor2 \comparator/C1598  ( .a(a[456]), .b(b[456]), .out(\comparator/N1133 )
         );
  xor2 \comparator/C1599  ( .a(a[455]), .b(b[455]), .out(\comparator/N1135 )
         );
  xor2 \comparator/C1600  ( .a(a[454]), .b(b[454]), .out(\comparator/N1137 )
         );
  xor2 \comparator/C1601  ( .a(a[453]), .b(b[453]), .out(\comparator/N1139 )
         );
  xor2 \comparator/C1602  ( .a(a[452]), .b(b[452]), .out(\comparator/N1141 )
         );
  xor2 \comparator/C1603  ( .a(a[451]), .b(b[451]), .out(\comparator/N1143 )
         );
  xor2 \comparator/C1604  ( .a(a[450]), .b(b[450]), .out(\comparator/N1145 )
         );
  xor2 \comparator/C1605  ( .a(a[449]), .b(b[449]), .out(\comparator/N1147 )
         );
  xor2 \comparator/C1606  ( .a(a[448]), .b(b[448]), .out(\comparator/N1149 )
         );
  xor2 \comparator/C1607  ( .a(a[447]), .b(b[447]), .out(\comparator/N1151 )
         );
  xor2 \comparator/C1608  ( .a(a[446]), .b(b[446]), .out(\comparator/N1153 )
         );
  xor2 \comparator/C1609  ( .a(a[445]), .b(b[445]), .out(\comparator/N1155 )
         );
  xor2 \comparator/C1610  ( .a(a[444]), .b(b[444]), .out(\comparator/N1157 )
         );
  xor2 \comparator/C1611  ( .a(a[443]), .b(b[443]), .out(\comparator/N1159 )
         );
  xor2 \comparator/C1612  ( .a(a[442]), .b(b[442]), .out(\comparator/N1161 )
         );
  xor2 \comparator/C1613  ( .a(a[441]), .b(b[441]), .out(\comparator/N1163 )
         );
  xor2 \comparator/C1614  ( .a(a[440]), .b(b[440]), .out(\comparator/N1165 )
         );
  xor2 \comparator/C1615  ( .a(a[439]), .b(b[439]), .out(\comparator/N1167 )
         );
  xor2 \comparator/C1616  ( .a(a[438]), .b(b[438]), .out(\comparator/N1169 )
         );
  xor2 \comparator/C1617  ( .a(a[437]), .b(b[437]), .out(\comparator/N1171 )
         );
  xor2 \comparator/C1618  ( .a(a[436]), .b(b[436]), .out(\comparator/N1173 )
         );
  xor2 \comparator/C1619  ( .a(a[435]), .b(b[435]), .out(\comparator/N1175 )
         );
  xor2 \comparator/C1620  ( .a(a[434]), .b(b[434]), .out(\comparator/N1177 )
         );
  xor2 \comparator/C1621  ( .a(a[433]), .b(b[433]), .out(\comparator/N1179 )
         );
  xor2 \comparator/C1622  ( .a(a[432]), .b(b[432]), .out(\comparator/N1181 )
         );
  xor2 \comparator/C1623  ( .a(a[431]), .b(b[431]), .out(\comparator/N1183 )
         );
  xor2 \comparator/C1624  ( .a(a[430]), .b(b[430]), .out(\comparator/N1185 )
         );
  xor2 \comparator/C1625  ( .a(a[429]), .b(b[429]), .out(\comparator/N1187 )
         );
  xor2 \comparator/C1626  ( .a(a[428]), .b(b[428]), .out(\comparator/N1189 )
         );
  xor2 \comparator/C1627  ( .a(a[427]), .b(b[427]), .out(\comparator/N1191 )
         );
  xor2 \comparator/C1628  ( .a(a[426]), .b(b[426]), .out(\comparator/N1193 )
         );
  xor2 \comparator/C1629  ( .a(a[425]), .b(b[425]), .out(\comparator/N1195 )
         );
  xor2 \comparator/C1630  ( .a(a[424]), .b(b[424]), .out(\comparator/N1197 )
         );
  xor2 \comparator/C1631  ( .a(a[423]), .b(b[423]), .out(\comparator/N1199 )
         );
  xor2 \comparator/C1632  ( .a(a[422]), .b(b[422]), .out(\comparator/N1201 )
         );
  xor2 \comparator/C1633  ( .a(a[421]), .b(b[421]), .out(\comparator/N1203 )
         );
  xor2 \comparator/C1634  ( .a(a[420]), .b(b[420]), .out(\comparator/N1205 )
         );
  xor2 \comparator/C1635  ( .a(a[419]), .b(b[419]), .out(\comparator/N1207 )
         );
  xor2 \comparator/C1636  ( .a(a[418]), .b(b[418]), .out(\comparator/N1209 )
         );
  xor2 \comparator/C1637  ( .a(a[417]), .b(b[417]), .out(\comparator/N1211 )
         );
  xor2 \comparator/C1638  ( .a(a[416]), .b(b[416]), .out(\comparator/N1213 )
         );
  xor2 \comparator/C1639  ( .a(a[415]), .b(b[415]), .out(\comparator/N1215 )
         );
  xor2 \comparator/C1640  ( .a(a[414]), .b(b[414]), .out(\comparator/N1217 )
         );
  xor2 \comparator/C1641  ( .a(a[413]), .b(b[413]), .out(\comparator/N1219 )
         );
  xor2 \comparator/C1642  ( .a(a[412]), .b(b[412]), .out(\comparator/N1221 )
         );
  xor2 \comparator/C1643  ( .a(a[411]), .b(b[411]), .out(\comparator/N1223 )
         );
  xor2 \comparator/C1644  ( .a(a[410]), .b(b[410]), .out(\comparator/N1225 )
         );
  xor2 \comparator/C1645  ( .a(a[409]), .b(b[409]), .out(\comparator/N1227 )
         );
  xor2 \comparator/C1646  ( .a(a[408]), .b(b[408]), .out(\comparator/N1229 )
         );
  xor2 \comparator/C1647  ( .a(a[407]), .b(b[407]), .out(\comparator/N1231 )
         );
  xor2 \comparator/C1648  ( .a(a[406]), .b(b[406]), .out(\comparator/N1233 )
         );
  xor2 \comparator/C1649  ( .a(a[405]), .b(b[405]), .out(\comparator/N1235 )
         );
  xor2 \comparator/C1650  ( .a(a[404]), .b(b[404]), .out(\comparator/N1237 )
         );
  xor2 \comparator/C1651  ( .a(a[403]), .b(b[403]), .out(\comparator/N1239 )
         );
  xor2 \comparator/C1652  ( .a(a[402]), .b(b[402]), .out(\comparator/N1241 )
         );
  xor2 \comparator/C1653  ( .a(a[401]), .b(b[401]), .out(\comparator/N1243 )
         );
  xor2 \comparator/C1654  ( .a(a[400]), .b(b[400]), .out(\comparator/N1245 )
         );
  xor2 \comparator/C1655  ( .a(a[399]), .b(b[399]), .out(\comparator/N1247 )
         );
  xor2 \comparator/C1656  ( .a(a[398]), .b(b[398]), .out(\comparator/N1249 )
         );
  xor2 \comparator/C1657  ( .a(a[397]), .b(b[397]), .out(\comparator/N1251 )
         );
  xor2 \comparator/C1658  ( .a(a[396]), .b(b[396]), .out(\comparator/N1253 )
         );
  xor2 \comparator/C1659  ( .a(a[395]), .b(b[395]), .out(\comparator/N1255 )
         );
  xor2 \comparator/C1660  ( .a(a[394]), .b(b[394]), .out(\comparator/N1257 )
         );
  xor2 \comparator/C1661  ( .a(a[393]), .b(b[393]), .out(\comparator/N1259 )
         );
  xor2 \comparator/C1662  ( .a(a[392]), .b(b[392]), .out(\comparator/N1261 )
         );
  xor2 \comparator/C1663  ( .a(a[391]), .b(b[391]), .out(\comparator/N1263 )
         );
  xor2 \comparator/C1664  ( .a(a[390]), .b(b[390]), .out(\comparator/N1265 )
         );
  xor2 \comparator/C1665  ( .a(a[389]), .b(b[389]), .out(\comparator/N1267 )
         );
  xor2 \comparator/C1666  ( .a(a[388]), .b(b[388]), .out(\comparator/N1269 )
         );
  xor2 \comparator/C1667  ( .a(a[387]), .b(b[387]), .out(\comparator/N1271 )
         );
  xor2 \comparator/C1668  ( .a(a[386]), .b(b[386]), .out(\comparator/N1273 )
         );
  xor2 \comparator/C1669  ( .a(a[385]), .b(b[385]), .out(\comparator/N1275 )
         );
  xor2 \comparator/C1670  ( .a(a[384]), .b(b[384]), .out(\comparator/N1277 )
         );
  xor2 \comparator/C1671  ( .a(a[383]), .b(b[383]), .out(\comparator/N1279 )
         );
  xor2 \comparator/C1672  ( .a(a[382]), .b(b[382]), .out(\comparator/N1281 )
         );
  xor2 \comparator/C1673  ( .a(a[381]), .b(b[381]), .out(\comparator/N1283 )
         );
  xor2 \comparator/C1674  ( .a(a[380]), .b(b[380]), .out(\comparator/N1285 )
         );
  xor2 \comparator/C1675  ( .a(a[379]), .b(b[379]), .out(\comparator/N1287 )
         );
  xor2 \comparator/C1676  ( .a(a[378]), .b(b[378]), .out(\comparator/N1289 )
         );
  xor2 \comparator/C1677  ( .a(a[377]), .b(b[377]), .out(\comparator/N1291 )
         );
  xor2 \comparator/C1678  ( .a(a[376]), .b(b[376]), .out(\comparator/N1293 )
         );
  xor2 \comparator/C1679  ( .a(a[375]), .b(b[375]), .out(\comparator/N1295 )
         );
  xor2 \comparator/C1680  ( .a(a[374]), .b(b[374]), .out(\comparator/N1297 )
         );
  xor2 \comparator/C1681  ( .a(a[373]), .b(b[373]), .out(\comparator/N1299 )
         );
  xor2 \comparator/C1682  ( .a(a[372]), .b(b[372]), .out(\comparator/N1301 )
         );
  xor2 \comparator/C1683  ( .a(a[371]), .b(b[371]), .out(\comparator/N1303 )
         );
  xor2 \comparator/C1684  ( .a(a[370]), .b(b[370]), .out(\comparator/N1305 )
         );
  xor2 \comparator/C1685  ( .a(a[369]), .b(b[369]), .out(\comparator/N1307 )
         );
  xor2 \comparator/C1686  ( .a(a[368]), .b(b[368]), .out(\comparator/N1309 )
         );
  xor2 \comparator/C1687  ( .a(a[367]), .b(b[367]), .out(\comparator/N1311 )
         );
  xor2 \comparator/C1688  ( .a(a[366]), .b(b[366]), .out(\comparator/N1313 )
         );
  xor2 \comparator/C1689  ( .a(a[365]), .b(b[365]), .out(\comparator/N1315 )
         );
  xor2 \comparator/C1690  ( .a(a[364]), .b(b[364]), .out(\comparator/N1317 )
         );
  xor2 \comparator/C1691  ( .a(a[363]), .b(b[363]), .out(\comparator/N1319 )
         );
  xor2 \comparator/C1692  ( .a(a[362]), .b(b[362]), .out(\comparator/N1321 )
         );
  xor2 \comparator/C1693  ( .a(a[361]), .b(b[361]), .out(\comparator/N1323 )
         );
  xor2 \comparator/C1694  ( .a(a[360]), .b(b[360]), .out(\comparator/N1325 )
         );
  xor2 \comparator/C1695  ( .a(a[359]), .b(b[359]), .out(\comparator/N1327 )
         );
  xor2 \comparator/C1696  ( .a(a[358]), .b(b[358]), .out(\comparator/N1329 )
         );
  xor2 \comparator/C1697  ( .a(a[357]), .b(b[357]), .out(\comparator/N1331 )
         );
  xor2 \comparator/C1698  ( .a(a[356]), .b(b[356]), .out(\comparator/N1333 )
         );
  xor2 \comparator/C1699  ( .a(a[355]), .b(b[355]), .out(\comparator/N1335 )
         );
  xor2 \comparator/C1700  ( .a(a[354]), .b(b[354]), .out(\comparator/N1337 )
         );
  xor2 \comparator/C1701  ( .a(a[353]), .b(b[353]), .out(\comparator/N1339 )
         );
  xor2 \comparator/C1702  ( .a(a[352]), .b(b[352]), .out(\comparator/N1341 )
         );
  xor2 \comparator/C1703  ( .a(a[351]), .b(b[351]), .out(\comparator/N1343 )
         );
  xor2 \comparator/C1704  ( .a(a[350]), .b(b[350]), .out(\comparator/N1345 )
         );
  xor2 \comparator/C1705  ( .a(a[349]), .b(b[349]), .out(\comparator/N1347 )
         );
  xor2 \comparator/C1706  ( .a(a[348]), .b(b[348]), .out(\comparator/N1349 )
         );
  xor2 \comparator/C1707  ( .a(a[347]), .b(b[347]), .out(\comparator/N1351 )
         );
  xor2 \comparator/C1708  ( .a(a[346]), .b(b[346]), .out(\comparator/N1353 )
         );
  xor2 \comparator/C1709  ( .a(a[345]), .b(b[345]), .out(\comparator/N1355 )
         );
  xor2 \comparator/C1710  ( .a(a[344]), .b(b[344]), .out(\comparator/N1357 )
         );
  xor2 \comparator/C1711  ( .a(a[343]), .b(b[343]), .out(\comparator/N1359 )
         );
  xor2 \comparator/C1712  ( .a(a[342]), .b(b[342]), .out(\comparator/N1361 )
         );
  xor2 \comparator/C1713  ( .a(a[341]), .b(b[341]), .out(\comparator/N1363 )
         );
  xor2 \comparator/C1714  ( .a(a[340]), .b(b[340]), .out(\comparator/N1365 )
         );
  xor2 \comparator/C1715  ( .a(a[339]), .b(b[339]), .out(\comparator/N1367 )
         );
  xor2 \comparator/C1716  ( .a(a[338]), .b(b[338]), .out(\comparator/N1369 )
         );
  xor2 \comparator/C1717  ( .a(a[337]), .b(b[337]), .out(\comparator/N1371 )
         );
  xor2 \comparator/C1718  ( .a(a[336]), .b(b[336]), .out(\comparator/N1373 )
         );
  xor2 \comparator/C1719  ( .a(a[335]), .b(b[335]), .out(\comparator/N1375 )
         );
  xor2 \comparator/C1720  ( .a(a[334]), .b(b[334]), .out(\comparator/N1377 )
         );
  xor2 \comparator/C1721  ( .a(a[333]), .b(b[333]), .out(\comparator/N1379 )
         );
  xor2 \comparator/C1722  ( .a(a[332]), .b(b[332]), .out(\comparator/N1381 )
         );
  xor2 \comparator/C1723  ( .a(a[331]), .b(b[331]), .out(\comparator/N1383 )
         );
  xor2 \comparator/C1724  ( .a(a[330]), .b(b[330]), .out(\comparator/N1385 )
         );
  xor2 \comparator/C1725  ( .a(a[329]), .b(b[329]), .out(\comparator/N1387 )
         );
  xor2 \comparator/C1726  ( .a(a[328]), .b(b[328]), .out(\comparator/N1389 )
         );
  xor2 \comparator/C1727  ( .a(a[327]), .b(b[327]), .out(\comparator/N1391 )
         );
  xor2 \comparator/C1728  ( .a(a[326]), .b(b[326]), .out(\comparator/N1393 )
         );
  xor2 \comparator/C1729  ( .a(a[325]), .b(b[325]), .out(\comparator/N1395 )
         );
  xor2 \comparator/C1730  ( .a(a[324]), .b(b[324]), .out(\comparator/N1397 )
         );
  xor2 \comparator/C1731  ( .a(a[323]), .b(b[323]), .out(\comparator/N1399 )
         );
  xor2 \comparator/C1732  ( .a(a[322]), .b(b[322]), .out(\comparator/N1401 )
         );
  xor2 \comparator/C1733  ( .a(a[321]), .b(b[321]), .out(\comparator/N1403 )
         );
  xor2 \comparator/C1734  ( .a(a[320]), .b(b[320]), .out(\comparator/N1405 )
         );
  xor2 \comparator/C1735  ( .a(a[319]), .b(b[319]), .out(\comparator/N1407 )
         );
  xor2 \comparator/C1736  ( .a(a[318]), .b(b[318]), .out(\comparator/N1409 )
         );
  xor2 \comparator/C1737  ( .a(a[317]), .b(b[317]), .out(\comparator/N1411 )
         );
  xor2 \comparator/C1738  ( .a(a[316]), .b(b[316]), .out(\comparator/N1413 )
         );
  xor2 \comparator/C1739  ( .a(a[315]), .b(b[315]), .out(\comparator/N1415 )
         );
  xor2 \comparator/C1740  ( .a(a[314]), .b(b[314]), .out(\comparator/N1417 )
         );
  xor2 \comparator/C1741  ( .a(a[313]), .b(b[313]), .out(\comparator/N1419 )
         );
  xor2 \comparator/C1742  ( .a(a[312]), .b(b[312]), .out(\comparator/N1421 )
         );
  xor2 \comparator/C1743  ( .a(a[311]), .b(b[311]), .out(\comparator/N1423 )
         );
  xor2 \comparator/C1744  ( .a(a[310]), .b(b[310]), .out(\comparator/N1425 )
         );
  xor2 \comparator/C1745  ( .a(a[309]), .b(b[309]), .out(\comparator/N1427 )
         );
  xor2 \comparator/C1746  ( .a(a[308]), .b(b[308]), .out(\comparator/N1429 )
         );
  xor2 \comparator/C1747  ( .a(a[307]), .b(b[307]), .out(\comparator/N1431 )
         );
  xor2 \comparator/C1748  ( .a(a[306]), .b(b[306]), .out(\comparator/N1433 )
         );
  xor2 \comparator/C1749  ( .a(a[305]), .b(b[305]), .out(\comparator/N1435 )
         );
  xor2 \comparator/C1750  ( .a(a[304]), .b(b[304]), .out(\comparator/N1437 )
         );
  xor2 \comparator/C1751  ( .a(a[303]), .b(b[303]), .out(\comparator/N1439 )
         );
  xor2 \comparator/C1752  ( .a(a[302]), .b(b[302]), .out(\comparator/N1441 )
         );
  xor2 \comparator/C1753  ( .a(a[301]), .b(b[301]), .out(\comparator/N1443 )
         );
  xor2 \comparator/C1754  ( .a(a[300]), .b(b[300]), .out(\comparator/N1445 )
         );
  xor2 \comparator/C1755  ( .a(a[299]), .b(b[299]), .out(\comparator/N1447 )
         );
  xor2 \comparator/C1756  ( .a(a[298]), .b(b[298]), .out(\comparator/N1449 )
         );
  xor2 \comparator/C1757  ( .a(a[297]), .b(b[297]), .out(\comparator/N1451 )
         );
  xor2 \comparator/C1758  ( .a(a[296]), .b(b[296]), .out(\comparator/N1453 )
         );
  xor2 \comparator/C1759  ( .a(a[295]), .b(b[295]), .out(\comparator/N1455 )
         );
  xor2 \comparator/C1760  ( .a(a[294]), .b(b[294]), .out(\comparator/N1457 )
         );
  xor2 \comparator/C1761  ( .a(a[293]), .b(b[293]), .out(\comparator/N1459 )
         );
  xor2 \comparator/C1762  ( .a(a[292]), .b(b[292]), .out(\comparator/N1461 )
         );
  xor2 \comparator/C1763  ( .a(a[291]), .b(b[291]), .out(\comparator/N1463 )
         );
  xor2 \comparator/C1764  ( .a(a[290]), .b(b[290]), .out(\comparator/N1465 )
         );
  xor2 \comparator/C1765  ( .a(a[289]), .b(b[289]), .out(\comparator/N1467 )
         );
  xor2 \comparator/C1766  ( .a(a[288]), .b(b[288]), .out(\comparator/N1469 )
         );
  xor2 \comparator/C1767  ( .a(a[287]), .b(b[287]), .out(\comparator/N1471 )
         );
  xor2 \comparator/C1768  ( .a(a[286]), .b(b[286]), .out(\comparator/N1473 )
         );
  xor2 \comparator/C1769  ( .a(a[285]), .b(b[285]), .out(\comparator/N1475 )
         );
  xor2 \comparator/C1770  ( .a(a[284]), .b(b[284]), .out(\comparator/N1477 )
         );
  xor2 \comparator/C1771  ( .a(a[283]), .b(b[283]), .out(\comparator/N1479 )
         );
  xor2 \comparator/C1772  ( .a(a[282]), .b(b[282]), .out(\comparator/N1481 )
         );
  xor2 \comparator/C1773  ( .a(a[281]), .b(b[281]), .out(\comparator/N1483 )
         );
  xor2 \comparator/C1774  ( .a(a[280]), .b(b[280]), .out(\comparator/N1485 )
         );
  xor2 \comparator/C1775  ( .a(a[279]), .b(b[279]), .out(\comparator/N1487 )
         );
  xor2 \comparator/C1776  ( .a(a[278]), .b(b[278]), .out(\comparator/N1489 )
         );
  xor2 \comparator/C1777  ( .a(a[277]), .b(b[277]), .out(\comparator/N1491 )
         );
  xor2 \comparator/C1778  ( .a(a[276]), .b(b[276]), .out(\comparator/N1493 )
         );
  xor2 \comparator/C1779  ( .a(a[275]), .b(b[275]), .out(\comparator/N1495 )
         );
  xor2 \comparator/C1780  ( .a(a[274]), .b(b[274]), .out(\comparator/N1497 )
         );
  xor2 \comparator/C1781  ( .a(a[273]), .b(b[273]), .out(\comparator/N1499 )
         );
  xor2 \comparator/C1782  ( .a(a[272]), .b(b[272]), .out(\comparator/N1501 )
         );
  xor2 \comparator/C1783  ( .a(a[271]), .b(b[271]), .out(\comparator/N1503 )
         );
  xor2 \comparator/C1784  ( .a(a[270]), .b(b[270]), .out(\comparator/N1505 )
         );
  xor2 \comparator/C1785  ( .a(a[269]), .b(b[269]), .out(\comparator/N1507 )
         );
  xor2 \comparator/C1786  ( .a(a[268]), .b(b[268]), .out(\comparator/N1509 )
         );
  xor2 \comparator/C1787  ( .a(a[267]), .b(b[267]), .out(\comparator/N1511 )
         );
  xor2 \comparator/C1788  ( .a(a[266]), .b(b[266]), .out(\comparator/N1513 )
         );
  xor2 \comparator/C1789  ( .a(a[265]), .b(b[265]), .out(\comparator/N1515 )
         );
  xor2 \comparator/C1790  ( .a(a[264]), .b(b[264]), .out(\comparator/N1517 )
         );
  xor2 \comparator/C1791  ( .a(a[263]), .b(b[263]), .out(\comparator/N1519 )
         );
  xor2 \comparator/C1792  ( .a(a[262]), .b(b[262]), .out(\comparator/N1521 )
         );
  xor2 \comparator/C1793  ( .a(a[261]), .b(b[261]), .out(\comparator/N1523 )
         );
  xor2 \comparator/C1794  ( .a(a[260]), .b(b[260]), .out(\comparator/N1525 )
         );
  xor2 \comparator/C1795  ( .a(a[259]), .b(b[259]), .out(\comparator/N1527 )
         );
  xor2 \comparator/C1796  ( .a(a[258]), .b(b[258]), .out(\comparator/N1529 )
         );
  xor2 \comparator/C1797  ( .a(a[257]), .b(b[257]), .out(\comparator/N1531 )
         );
  xor2 \comparator/C1798  ( .a(a[256]), .b(b[256]), .out(\comparator/N1533 )
         );
  xor2 \comparator/C1799  ( .a(a[255]), .b(b[255]), .out(\comparator/N1535 )
         );
  xor2 \comparator/C1800  ( .a(a[254]), .b(b[254]), .out(\comparator/N1537 )
         );
  xor2 \comparator/C1801  ( .a(a[253]), .b(b[253]), .out(\comparator/N1539 )
         );
  xor2 \comparator/C1802  ( .a(a[252]), .b(b[252]), .out(\comparator/N1541 )
         );
  xor2 \comparator/C1803  ( .a(a[251]), .b(b[251]), .out(\comparator/N1543 )
         );
  xor2 \comparator/C1804  ( .a(a[250]), .b(b[250]), .out(\comparator/N1545 )
         );
  xor2 \comparator/C1805  ( .a(a[249]), .b(b[249]), .out(\comparator/N1547 )
         );
  xor2 \comparator/C1806  ( .a(a[248]), .b(b[248]), .out(\comparator/N1549 )
         );
  xor2 \comparator/C1807  ( .a(a[247]), .b(b[247]), .out(\comparator/N1551 )
         );
  xor2 \comparator/C1808  ( .a(a[246]), .b(b[246]), .out(\comparator/N1553 )
         );
  xor2 \comparator/C1809  ( .a(a[245]), .b(b[245]), .out(\comparator/N1555 )
         );
  xor2 \comparator/C1810  ( .a(a[244]), .b(b[244]), .out(\comparator/N1557 )
         );
  xor2 \comparator/C1811  ( .a(a[243]), .b(b[243]), .out(\comparator/N1559 )
         );
  xor2 \comparator/C1812  ( .a(a[242]), .b(b[242]), .out(\comparator/N1561 )
         );
  xor2 \comparator/C1813  ( .a(a[241]), .b(b[241]), .out(\comparator/N1563 )
         );
  xor2 \comparator/C1814  ( .a(a[240]), .b(b[240]), .out(\comparator/N1565 )
         );
  xor2 \comparator/C1815  ( .a(a[239]), .b(b[239]), .out(\comparator/N1567 )
         );
  xor2 \comparator/C1816  ( .a(a[238]), .b(b[238]), .out(\comparator/N1569 )
         );
  xor2 \comparator/C1817  ( .a(a[237]), .b(b[237]), .out(\comparator/N1571 )
         );
  xor2 \comparator/C1818  ( .a(a[236]), .b(b[236]), .out(\comparator/N1573 )
         );
  xor2 \comparator/C1819  ( .a(a[235]), .b(b[235]), .out(\comparator/N1575 )
         );
  xor2 \comparator/C1820  ( .a(a[234]), .b(b[234]), .out(\comparator/N1577 )
         );
  xor2 \comparator/C1821  ( .a(a[233]), .b(b[233]), .out(\comparator/N1579 )
         );
  xor2 \comparator/C1822  ( .a(a[232]), .b(b[232]), .out(\comparator/N1581 )
         );
  xor2 \comparator/C1823  ( .a(a[231]), .b(b[231]), .out(\comparator/N1583 )
         );
  xor2 \comparator/C1824  ( .a(a[230]), .b(b[230]), .out(\comparator/N1585 )
         );
  xor2 \comparator/C1825  ( .a(a[229]), .b(b[229]), .out(\comparator/N1587 )
         );
  xor2 \comparator/C1826  ( .a(a[228]), .b(b[228]), .out(\comparator/N1589 )
         );
  xor2 \comparator/C1827  ( .a(a[227]), .b(b[227]), .out(\comparator/N1591 )
         );
  xor2 \comparator/C1828  ( .a(a[226]), .b(b[226]), .out(\comparator/N1593 )
         );
  xor2 \comparator/C1829  ( .a(a[225]), .b(b[225]), .out(\comparator/N1595 )
         );
  xor2 \comparator/C1830  ( .a(a[224]), .b(b[224]), .out(\comparator/N1597 )
         );
  xor2 \comparator/C1831  ( .a(a[223]), .b(b[223]), .out(\comparator/N1599 )
         );
  xor2 \comparator/C1832  ( .a(a[222]), .b(b[222]), .out(\comparator/N1601 )
         );
  xor2 \comparator/C1833  ( .a(a[221]), .b(b[221]), .out(\comparator/N1603 )
         );
  xor2 \comparator/C1834  ( .a(a[220]), .b(b[220]), .out(\comparator/N1605 )
         );
  xor2 \comparator/C1835  ( .a(a[219]), .b(b[219]), .out(\comparator/N1607 )
         );
  xor2 \comparator/C1836  ( .a(a[218]), .b(b[218]), .out(\comparator/N1609 )
         );
  xor2 \comparator/C1837  ( .a(a[217]), .b(b[217]), .out(\comparator/N1611 )
         );
  xor2 \comparator/C1838  ( .a(a[216]), .b(b[216]), .out(\comparator/N1613 )
         );
  xor2 \comparator/C1839  ( .a(a[215]), .b(b[215]), .out(\comparator/N1615 )
         );
  xor2 \comparator/C1840  ( .a(a[214]), .b(b[214]), .out(\comparator/N1617 )
         );
  xor2 \comparator/C1841  ( .a(a[213]), .b(b[213]), .out(\comparator/N1619 )
         );
  xor2 \comparator/C1842  ( .a(a[212]), .b(b[212]), .out(\comparator/N1621 )
         );
  xor2 \comparator/C1843  ( .a(a[211]), .b(b[211]), .out(\comparator/N1623 )
         );
  xor2 \comparator/C1844  ( .a(a[210]), .b(b[210]), .out(\comparator/N1625 )
         );
  xor2 \comparator/C1845  ( .a(a[209]), .b(b[209]), .out(\comparator/N1627 )
         );
  xor2 \comparator/C1846  ( .a(a[208]), .b(b[208]), .out(\comparator/N1629 )
         );
  xor2 \comparator/C1847  ( .a(a[207]), .b(b[207]), .out(\comparator/N1631 )
         );
  xor2 \comparator/C1848  ( .a(a[206]), .b(b[206]), .out(\comparator/N1633 )
         );
  xor2 \comparator/C1849  ( .a(a[205]), .b(b[205]), .out(\comparator/N1635 )
         );
  xor2 \comparator/C1850  ( .a(a[204]), .b(b[204]), .out(\comparator/N1637 )
         );
  xor2 \comparator/C1851  ( .a(a[203]), .b(b[203]), .out(\comparator/N1639 )
         );
  xor2 \comparator/C1852  ( .a(a[202]), .b(b[202]), .out(\comparator/N1641 )
         );
  xor2 \comparator/C1853  ( .a(a[201]), .b(b[201]), .out(\comparator/N1643 )
         );
  xor2 \comparator/C1854  ( .a(a[200]), .b(b[200]), .out(\comparator/N1645 )
         );
  xor2 \comparator/C1855  ( .a(a[199]), .b(b[199]), .out(\comparator/N1647 )
         );
  xor2 \comparator/C1856  ( .a(a[198]), .b(b[198]), .out(\comparator/N1649 )
         );
  xor2 \comparator/C1857  ( .a(a[197]), .b(b[197]), .out(\comparator/N1651 )
         );
  xor2 \comparator/C1858  ( .a(a[196]), .b(b[196]), .out(\comparator/N1653 )
         );
  xor2 \comparator/C1859  ( .a(a[195]), .b(b[195]), .out(\comparator/N1655 )
         );
  xor2 \comparator/C1860  ( .a(a[194]), .b(b[194]), .out(\comparator/N1657 )
         );
  xor2 \comparator/C1861  ( .a(a[193]), .b(b[193]), .out(\comparator/N1659 )
         );
  xor2 \comparator/C1862  ( .a(a[192]), .b(b[192]), .out(\comparator/N1661 )
         );
  xor2 \comparator/C1863  ( .a(a[191]), .b(b[191]), .out(\comparator/N1663 )
         );
  xor2 \comparator/C1864  ( .a(a[190]), .b(b[190]), .out(\comparator/N1665 )
         );
  xor2 \comparator/C1865  ( .a(a[189]), .b(b[189]), .out(\comparator/N1667 )
         );
  xor2 \comparator/C1866  ( .a(a[188]), .b(b[188]), .out(\comparator/N1669 )
         );
  xor2 \comparator/C1867  ( .a(a[187]), .b(b[187]), .out(\comparator/N1671 )
         );
  xor2 \comparator/C1868  ( .a(a[186]), .b(b[186]), .out(\comparator/N1673 )
         );
  xor2 \comparator/C1869  ( .a(a[185]), .b(b[185]), .out(\comparator/N1675 )
         );
  xor2 \comparator/C1870  ( .a(a[184]), .b(b[184]), .out(\comparator/N1677 )
         );
  xor2 \comparator/C1871  ( .a(a[183]), .b(b[183]), .out(\comparator/N1679 )
         );
  xor2 \comparator/C1872  ( .a(a[182]), .b(b[182]), .out(\comparator/N1681 )
         );
  xor2 \comparator/C1873  ( .a(a[181]), .b(b[181]), .out(\comparator/N1683 )
         );
  xor2 \comparator/C1874  ( .a(a[180]), .b(b[180]), .out(\comparator/N1685 )
         );
  xor2 \comparator/C1875  ( .a(a[179]), .b(b[179]), .out(\comparator/N1687 )
         );
  xor2 \comparator/C1876  ( .a(a[178]), .b(b[178]), .out(\comparator/N1689 )
         );
  xor2 \comparator/C1877  ( .a(a[177]), .b(b[177]), .out(\comparator/N1691 )
         );
  xor2 \comparator/C1878  ( .a(a[176]), .b(b[176]), .out(\comparator/N1693 )
         );
  xor2 \comparator/C1879  ( .a(a[175]), .b(b[175]), .out(\comparator/N1695 )
         );
  xor2 \comparator/C1880  ( .a(a[174]), .b(b[174]), .out(\comparator/N1697 )
         );
  xor2 \comparator/C1881  ( .a(a[173]), .b(b[173]), .out(\comparator/N1699 )
         );
  xor2 \comparator/C1882  ( .a(a[172]), .b(b[172]), .out(\comparator/N1701 )
         );
  xor2 \comparator/C1883  ( .a(a[171]), .b(b[171]), .out(\comparator/N1703 )
         );
  xor2 \comparator/C1884  ( .a(a[170]), .b(b[170]), .out(\comparator/N1705 )
         );
  xor2 \comparator/C1885  ( .a(a[169]), .b(b[169]), .out(\comparator/N1707 )
         );
  xor2 \comparator/C1886  ( .a(a[168]), .b(b[168]), .out(\comparator/N1709 )
         );
  xor2 \comparator/C1887  ( .a(a[167]), .b(b[167]), .out(\comparator/N1711 )
         );
  xor2 \comparator/C1888  ( .a(a[166]), .b(b[166]), .out(\comparator/N1713 )
         );
  xor2 \comparator/C1889  ( .a(a[165]), .b(b[165]), .out(\comparator/N1715 )
         );
  xor2 \comparator/C1890  ( .a(a[164]), .b(b[164]), .out(\comparator/N1717 )
         );
  xor2 \comparator/C1891  ( .a(a[163]), .b(b[163]), .out(\comparator/N1719 )
         );
  xor2 \comparator/C1892  ( .a(a[162]), .b(b[162]), .out(\comparator/N1721 )
         );
  xor2 \comparator/C1893  ( .a(a[161]), .b(b[161]), .out(\comparator/N1723 )
         );
  xor2 \comparator/C1894  ( .a(a[160]), .b(b[160]), .out(\comparator/N1725 )
         );
  xor2 \comparator/C1895  ( .a(a[159]), .b(b[159]), .out(\comparator/N1727 )
         );
  xor2 \comparator/C1896  ( .a(a[158]), .b(b[158]), .out(\comparator/N1729 )
         );
  xor2 \comparator/C1897  ( .a(a[157]), .b(b[157]), .out(\comparator/N1731 )
         );
  xor2 \comparator/C1898  ( .a(a[156]), .b(b[156]), .out(\comparator/N1733 )
         );
  xor2 \comparator/C1899  ( .a(a[155]), .b(b[155]), .out(\comparator/N1735 )
         );
  xor2 \comparator/C1900  ( .a(a[154]), .b(b[154]), .out(\comparator/N1737 )
         );
  xor2 \comparator/C1901  ( .a(a[153]), .b(b[153]), .out(\comparator/N1739 )
         );
  xor2 \comparator/C1902  ( .a(a[152]), .b(b[152]), .out(\comparator/N1741 )
         );
  xor2 \comparator/C1903  ( .a(a[151]), .b(b[151]), .out(\comparator/N1743 )
         );
  xor2 \comparator/C1904  ( .a(a[150]), .b(b[150]), .out(\comparator/N1745 )
         );
  xor2 \comparator/C1905  ( .a(a[149]), .b(b[149]), .out(\comparator/N1747 )
         );
  xor2 \comparator/C1906  ( .a(a[148]), .b(b[148]), .out(\comparator/N1749 )
         );
  xor2 \comparator/C1907  ( .a(a[147]), .b(b[147]), .out(\comparator/N1751 )
         );
  xor2 \comparator/C1908  ( .a(a[146]), .b(b[146]), .out(\comparator/N1753 )
         );
  xor2 \comparator/C1909  ( .a(a[145]), .b(b[145]), .out(\comparator/N1755 )
         );
  xor2 \comparator/C1910  ( .a(a[144]), .b(b[144]), .out(\comparator/N1757 )
         );
  xor2 \comparator/C1911  ( .a(a[143]), .b(b[143]), .out(\comparator/N1759 )
         );
  xor2 \comparator/C1912  ( .a(a[142]), .b(b[142]), .out(\comparator/N1761 )
         );
  xor2 \comparator/C1913  ( .a(a[141]), .b(b[141]), .out(\comparator/N1763 )
         );
  xor2 \comparator/C1914  ( .a(a[140]), .b(b[140]), .out(\comparator/N1765 )
         );
  xor2 \comparator/C1915  ( .a(a[139]), .b(b[139]), .out(\comparator/N1767 )
         );
  xor2 \comparator/C1916  ( .a(a[138]), .b(b[138]), .out(\comparator/N1769 )
         );
  xor2 \comparator/C1917  ( .a(a[137]), .b(b[137]), .out(\comparator/N1771 )
         );
  xor2 \comparator/C1918  ( .a(a[136]), .b(b[136]), .out(\comparator/N1773 )
         );
  xor2 \comparator/C1919  ( .a(a[135]), .b(b[135]), .out(\comparator/N1775 )
         );
  xor2 \comparator/C1920  ( .a(a[134]), .b(b[134]), .out(\comparator/N1777 )
         );
  xor2 \comparator/C1921  ( .a(a[133]), .b(b[133]), .out(\comparator/N1779 )
         );
  xor2 \comparator/C1922  ( .a(a[132]), .b(b[132]), .out(\comparator/N1781 )
         );
  xor2 \comparator/C1923  ( .a(a[131]), .b(b[131]), .out(\comparator/N1783 )
         );
  xor2 \comparator/C1924  ( .a(a[130]), .b(b[130]), .out(\comparator/N1785 )
         );
  xor2 \comparator/C1925  ( .a(a[129]), .b(b[129]), .out(\comparator/N1787 )
         );
  xor2 \comparator/C1926  ( .a(a[128]), .b(b[128]), .out(\comparator/N1789 )
         );
  xor2 \comparator/C1927  ( .a(a[127]), .b(b[127]), .out(\comparator/N1791 )
         );
  xor2 \comparator/C1928  ( .a(a[126]), .b(b[126]), .out(\comparator/N1793 )
         );
  xor2 \comparator/C1929  ( .a(a[125]), .b(b[125]), .out(\comparator/N1795 )
         );
  xor2 \comparator/C1930  ( .a(a[124]), .b(b[124]), .out(\comparator/N1797 )
         );
  xor2 \comparator/C1931  ( .a(a[123]), .b(b[123]), .out(\comparator/N1799 )
         );
  xor2 \comparator/C1932  ( .a(a[122]), .b(b[122]), .out(\comparator/N1801 )
         );
  xor2 \comparator/C1933  ( .a(a[121]), .b(b[121]), .out(\comparator/N1803 )
         );
  xor2 \comparator/C1934  ( .a(a[120]), .b(b[120]), .out(\comparator/N1805 )
         );
  xor2 \comparator/C1935  ( .a(a[119]), .b(b[119]), .out(\comparator/N1807 )
         );
  xor2 \comparator/C1936  ( .a(a[118]), .b(b[118]), .out(\comparator/N1809 )
         );
  xor2 \comparator/C1937  ( .a(a[117]), .b(b[117]), .out(\comparator/N1811 )
         );
  xor2 \comparator/C1938  ( .a(a[116]), .b(b[116]), .out(\comparator/N1813 )
         );
  xor2 \comparator/C1939  ( .a(a[115]), .b(b[115]), .out(\comparator/N1815 )
         );
  xor2 \comparator/C1940  ( .a(a[114]), .b(b[114]), .out(\comparator/N1817 )
         );
  xor2 \comparator/C1941  ( .a(a[113]), .b(b[113]), .out(\comparator/N1819 )
         );
  xor2 \comparator/C1942  ( .a(a[112]), .b(b[112]), .out(\comparator/N1821 )
         );
  xor2 \comparator/C1943  ( .a(a[111]), .b(b[111]), .out(\comparator/N1823 )
         );
  xor2 \comparator/C1944  ( .a(a[110]), .b(b[110]), .out(\comparator/N1825 )
         );
  xor2 \comparator/C1945  ( .a(a[109]), .b(b[109]), .out(\comparator/N1827 )
         );
  xor2 \comparator/C1946  ( .a(a[108]), .b(b[108]), .out(\comparator/N1829 )
         );
  xor2 \comparator/C1947  ( .a(a[107]), .b(b[107]), .out(\comparator/N1831 )
         );
  xor2 \comparator/C1948  ( .a(a[106]), .b(b[106]), .out(\comparator/N1833 )
         );
  xor2 \comparator/C1949  ( .a(a[105]), .b(b[105]), .out(\comparator/N1835 )
         );
  xor2 \comparator/C1950  ( .a(a[104]), .b(b[104]), .out(\comparator/N1837 )
         );
  xor2 \comparator/C1951  ( .a(a[103]), .b(b[103]), .out(\comparator/N1839 )
         );
  xor2 \comparator/C1952  ( .a(a[102]), .b(b[102]), .out(\comparator/N1841 )
         );
  xor2 \comparator/C1953  ( .a(a[101]), .b(b[101]), .out(\comparator/N1843 )
         );
  xor2 \comparator/C1954  ( .a(a[100]), .b(b[100]), .out(\comparator/N1845 )
         );
  xor2 \comparator/C1955  ( .a(a[99]), .b(b[99]), .out(\comparator/N1847 ) );
  xor2 \comparator/C1956  ( .a(a[98]), .b(b[98]), .out(\comparator/N1849 ) );
  xor2 \comparator/C1957  ( .a(a[97]), .b(b[97]), .out(\comparator/N1851 ) );
  xor2 \comparator/C1958  ( .a(a[96]), .b(b[96]), .out(\comparator/N1853 ) );
  xor2 \comparator/C1959  ( .a(a[95]), .b(b[95]), .out(\comparator/N1855 ) );
  xor2 \comparator/C1960  ( .a(a[94]), .b(b[94]), .out(\comparator/N1857 ) );
  xor2 \comparator/C1961  ( .a(a[93]), .b(b[93]), .out(\comparator/N1859 ) );
  xor2 \comparator/C1962  ( .a(a[92]), .b(b[92]), .out(\comparator/N1861 ) );
  xor2 \comparator/C1963  ( .a(a[91]), .b(b[91]), .out(\comparator/N1863 ) );
  xor2 \comparator/C1964  ( .a(a[90]), .b(b[90]), .out(\comparator/N1865 ) );
  xor2 \comparator/C1965  ( .a(a[89]), .b(b[89]), .out(\comparator/N1867 ) );
  xor2 \comparator/C1966  ( .a(a[88]), .b(b[88]), .out(\comparator/N1869 ) );
  xor2 \comparator/C1967  ( .a(a[87]), .b(b[87]), .out(\comparator/N1871 ) );
  xor2 \comparator/C1968  ( .a(a[86]), .b(b[86]), .out(\comparator/N1873 ) );
  xor2 \comparator/C1969  ( .a(a[85]), .b(b[85]), .out(\comparator/N1875 ) );
  xor2 \comparator/C1970  ( .a(a[84]), .b(b[84]), .out(\comparator/N1877 ) );
  xor2 \comparator/C1971  ( .a(a[83]), .b(b[83]), .out(\comparator/N1879 ) );
  xor2 \comparator/C1972  ( .a(a[82]), .b(b[82]), .out(\comparator/N1881 ) );
  xor2 \comparator/C1973  ( .a(a[81]), .b(b[81]), .out(\comparator/N1883 ) );
  xor2 \comparator/C1974  ( .a(a[80]), .b(b[80]), .out(\comparator/N1885 ) );
  xor2 \comparator/C1975  ( .a(a[79]), .b(b[79]), .out(\comparator/N1887 ) );
  xor2 \comparator/C1976  ( .a(a[78]), .b(b[78]), .out(\comparator/N1889 ) );
  xor2 \comparator/C1977  ( .a(a[77]), .b(b[77]), .out(\comparator/N1891 ) );
  xor2 \comparator/C1978  ( .a(a[76]), .b(b[76]), .out(\comparator/N1893 ) );
  xor2 \comparator/C1979  ( .a(a[75]), .b(b[75]), .out(\comparator/N1895 ) );
  xor2 \comparator/C1980  ( .a(a[74]), .b(b[74]), .out(\comparator/N1897 ) );
  xor2 \comparator/C1981  ( .a(a[73]), .b(b[73]), .out(\comparator/N1899 ) );
  xor2 \comparator/C1982  ( .a(a[72]), .b(b[72]), .out(\comparator/N1901 ) );
  xor2 \comparator/C1983  ( .a(a[71]), .b(b[71]), .out(\comparator/N1903 ) );
  xor2 \comparator/C1984  ( .a(a[70]), .b(b[70]), .out(\comparator/N1905 ) );
  xor2 \comparator/C1985  ( .a(a[69]), .b(b[69]), .out(\comparator/N1907 ) );
  xor2 \comparator/C1986  ( .a(a[68]), .b(b[68]), .out(\comparator/N1909 ) );
  xor2 \comparator/C1987  ( .a(a[67]), .b(b[67]), .out(\comparator/N1911 ) );
  xor2 \comparator/C1988  ( .a(a[66]), .b(b[66]), .out(\comparator/N1913 ) );
  xor2 \comparator/C1989  ( .a(a[65]), .b(b[65]), .out(\comparator/N1915 ) );
  xor2 \comparator/C1990  ( .a(a[64]), .b(b[64]), .out(\comparator/N1917 ) );
  xor2 \comparator/C1991  ( .a(a[63]), .b(b[63]), .out(\comparator/N1919 ) );
  xor2 \comparator/C1992  ( .a(a[62]), .b(b[62]), .out(\comparator/N1921 ) );
  xor2 \comparator/C1993  ( .a(a[61]), .b(b[61]), .out(\comparator/N1923 ) );
  xor2 \comparator/C1994  ( .a(a[60]), .b(b[60]), .out(\comparator/N1925 ) );
  xor2 \comparator/C1995  ( .a(a[59]), .b(b[59]), .out(\comparator/N1927 ) );
  xor2 \comparator/C1996  ( .a(a[58]), .b(b[58]), .out(\comparator/N1929 ) );
  xor2 \comparator/C1997  ( .a(a[57]), .b(b[57]), .out(\comparator/N1931 ) );
  xor2 \comparator/C1998  ( .a(a[56]), .b(b[56]), .out(\comparator/N1933 ) );
  xor2 \comparator/C1999  ( .a(a[55]), .b(b[55]), .out(\comparator/N1935 ) );
  xor2 \comparator/C2000  ( .a(a[54]), .b(b[54]), .out(\comparator/N1937 ) );
  xor2 \comparator/C2001  ( .a(a[53]), .b(b[53]), .out(\comparator/N1939 ) );
  xor2 \comparator/C2002  ( .a(a[52]), .b(b[52]), .out(\comparator/N1941 ) );
  xor2 \comparator/C2003  ( .a(a[51]), .b(b[51]), .out(\comparator/N1943 ) );
  xor2 \comparator/C2004  ( .a(a[50]), .b(b[50]), .out(\comparator/N1945 ) );
  xor2 \comparator/C2005  ( .a(a[49]), .b(b[49]), .out(\comparator/N1947 ) );
  xor2 \comparator/C2006  ( .a(a[48]), .b(b[48]), .out(\comparator/N1949 ) );
  xor2 \comparator/C2007  ( .a(a[47]), .b(b[47]), .out(\comparator/N1951 ) );
  xor2 \comparator/C2008  ( .a(a[46]), .b(b[46]), .out(\comparator/N1953 ) );
  xor2 \comparator/C2009  ( .a(a[45]), .b(b[45]), .out(\comparator/N1955 ) );
  xor2 \comparator/C2010  ( .a(a[44]), .b(b[44]), .out(\comparator/N1957 ) );
  xor2 \comparator/C2011  ( .a(a[43]), .b(b[43]), .out(\comparator/N1959 ) );
  xor2 \comparator/C2012  ( .a(a[42]), .b(b[42]), .out(\comparator/N1961 ) );
  xor2 \comparator/C2013  ( .a(a[41]), .b(b[41]), .out(\comparator/N1963 ) );
  xor2 \comparator/C2014  ( .a(a[40]), .b(b[40]), .out(\comparator/N1965 ) );
  xor2 \comparator/C2015  ( .a(a[39]), .b(b[39]), .out(\comparator/N1967 ) );
  xor2 \comparator/C2016  ( .a(a[38]), .b(b[38]), .out(\comparator/N1969 ) );
  xor2 \comparator/C2017  ( .a(a[37]), .b(b[37]), .out(\comparator/N1971 ) );
  xor2 \comparator/C2018  ( .a(a[36]), .b(b[36]), .out(\comparator/N1973 ) );
  xor2 \comparator/C2019  ( .a(a[35]), .b(b[35]), .out(\comparator/N1975 ) );
  xor2 \comparator/C2020  ( .a(a[34]), .b(b[34]), .out(\comparator/N1977 ) );
  xor2 \comparator/C2021  ( .a(a[33]), .b(b[33]), .out(\comparator/N1979 ) );
  xor2 \comparator/C2022  ( .a(a[32]), .b(b[32]), .out(\comparator/N1981 ) );
  xor2 \comparator/C2023  ( .a(a[31]), .b(b[31]), .out(\comparator/N1983 ) );
  xor2 \comparator/C2024  ( .a(a[30]), .b(b[30]), .out(\comparator/N1985 ) );
  xor2 \comparator/C2025  ( .a(a[29]), .b(b[29]), .out(\comparator/N1987 ) );
  xor2 \comparator/C2026  ( .a(a[28]), .b(b[28]), .out(\comparator/N1989 ) );
  xor2 \comparator/C2027  ( .a(a[27]), .b(b[27]), .out(\comparator/N1991 ) );
  xor2 \comparator/C2028  ( .a(a[26]), .b(b[26]), .out(\comparator/N1993 ) );
  xor2 \comparator/C2029  ( .a(a[25]), .b(b[25]), .out(\comparator/N1995 ) );
  xor2 \comparator/C2030  ( .a(a[24]), .b(b[24]), .out(\comparator/N1997 ) );
  xor2 \comparator/C2031  ( .a(a[23]), .b(b[23]), .out(\comparator/N1999 ) );
  xor2 \comparator/C2032  ( .a(a[22]), .b(b[22]), .out(\comparator/N2001 ) );
  xor2 \comparator/C2033  ( .a(a[21]), .b(b[21]), .out(\comparator/N2003 ) );
  xor2 \comparator/C2034  ( .a(a[20]), .b(b[20]), .out(\comparator/N2005 ) );
  xor2 \comparator/C2035  ( .a(a[19]), .b(b[19]), .out(\comparator/N2007 ) );
  xor2 \comparator/C2036  ( .a(a[18]), .b(b[18]), .out(\comparator/N2009 ) );
  xor2 \comparator/C2037  ( .a(a[17]), .b(b[17]), .out(\comparator/N2011 ) );
  xor2 \comparator/C2038  ( .a(a[16]), .b(b[16]), .out(\comparator/N2013 ) );
  xor2 \comparator/C2039  ( .a(a[15]), .b(b[15]), .out(\comparator/N2015 ) );
  xor2 \comparator/C2040  ( .a(a[14]), .b(b[14]), .out(\comparator/N2017 ) );
  xor2 \comparator/C2041  ( .a(a[13]), .b(b[13]), .out(\comparator/N2019 ) );
  xor2 \comparator/C2042  ( .a(a[12]), .b(b[12]), .out(\comparator/N2021 ) );
  xor2 \comparator/C2043  ( .a(a[11]), .b(b[11]), .out(\comparator/N2023 ) );
  xor2 \comparator/C2044  ( .a(a[10]), .b(b[10]), .out(\comparator/N2025 ) );
  xor2 \comparator/C2045  ( .a(a[9]), .b(b[9]), .out(\comparator/N2027 ) );
  xor2 \comparator/C2046  ( .a(a[8]), .b(b[8]), .out(\comparator/N2029 ) );
  xor2 \comparator/C2047  ( .a(a[7]), .b(b[7]), .out(\comparator/N2031 ) );
  xor2 \comparator/C2048  ( .a(a[6]), .b(b[6]), .out(\comparator/N2033 ) );
  xor2 \comparator/C2049  ( .a(a[5]), .b(b[5]), .out(\comparator/N2035 ) );
  xor2 \comparator/C2050  ( .a(a[4]), .b(b[4]), .out(\comparator/N2037 ) );
  xor2 \comparator/C2051  ( .a(a[3]), .b(b[3]), .out(\comparator/N2039 ) );
  xor2 \comparator/C2052  ( .a(a[2]), .b(b[2]), .out(\comparator/N2041 ) );
  xor2 \comparator/C2053  ( .a(a[1]), .b(b[1]), .out(\comparator/N2043 ) );
  xor2 \comparator/C2054  ( .a(a[0]), .b(b[0]), .out(\comparator/N2045 ) );
  inv \sig_prgm_register/I_0  ( .a(clr), .out(\sig_prgm_register/clear_not )
         );
  d_ff \sig_prgm_register/genblk1[1023].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1023]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1023]) );
  d_ff \sig_prgm_register/genblk1[1022].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1022]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1022]) );
  d_ff \sig_prgm_register/genblk1[1021].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1021]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1021]) );
  d_ff \sig_prgm_register/genblk1[1020].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1020]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1020]) );
  d_ff \sig_prgm_register/genblk1[1019].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1019]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1019]) );
  d_ff \sig_prgm_register/genblk1[1018].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1018]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1018]) );
  d_ff \sig_prgm_register/genblk1[1017].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1017]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1017]) );
  d_ff \sig_prgm_register/genblk1[1016].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1016]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1016]) );
  d_ff \sig_prgm_register/genblk1[1015].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1015]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1015]) );
  d_ff \sig_prgm_register/genblk1[1014].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1014]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1014]) );
  d_ff \sig_prgm_register/genblk1[1013].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1013]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1013]) );
  d_ff \sig_prgm_register/genblk1[1012].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1012]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1012]) );
  d_ff \sig_prgm_register/genblk1[1011].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1011]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1011]) );
  d_ff \sig_prgm_register/genblk1[1010].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1010]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1010]) );
  d_ff \sig_prgm_register/genblk1[1009].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1009]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1009]) );
  d_ff \sig_prgm_register/genblk1[1008].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1008]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1008]) );
  d_ff \sig_prgm_register/genblk1[1007].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1007]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1007]) );
  d_ff \sig_prgm_register/genblk1[1006].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1006]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1006]) );
  d_ff \sig_prgm_register/genblk1[1005].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1005]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1005]) );
  d_ff \sig_prgm_register/genblk1[1004].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1004]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1004]) );
  d_ff \sig_prgm_register/genblk1[1003].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1003]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1003]) );
  d_ff \sig_prgm_register/genblk1[1002].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1002]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1002]) );
  d_ff \sig_prgm_register/genblk1[1001].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1001]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1001]) );
  d_ff \sig_prgm_register/genblk1[1000].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1000]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1000]) );
  d_ff \sig_prgm_register/genblk1[999].single_DFF  ( .d(
        \sig_prgm_register/or_signal [999]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[999]) );
  d_ff \sig_prgm_register/genblk1[998].single_DFF  ( .d(
        \sig_prgm_register/or_signal [998]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[998]) );
  d_ff \sig_prgm_register/genblk1[997].single_DFF  ( .d(
        \sig_prgm_register/or_signal [997]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[997]) );
  d_ff \sig_prgm_register/genblk1[996].single_DFF  ( .d(
        \sig_prgm_register/or_signal [996]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[996]) );
  d_ff \sig_prgm_register/genblk1[995].single_DFF  ( .d(
        \sig_prgm_register/or_signal [995]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[995]) );
  d_ff \sig_prgm_register/genblk1[994].single_DFF  ( .d(
        \sig_prgm_register/or_signal [994]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[994]) );
  d_ff \sig_prgm_register/genblk1[993].single_DFF  ( .d(
        \sig_prgm_register/or_signal [993]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[993]) );
  d_ff \sig_prgm_register/genblk1[992].single_DFF  ( .d(
        \sig_prgm_register/or_signal [992]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[992]) );
  d_ff \sig_prgm_register/genblk1[991].single_DFF  ( .d(
        \sig_prgm_register/or_signal [991]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[991]) );
  d_ff \sig_prgm_register/genblk1[990].single_DFF  ( .d(
        \sig_prgm_register/or_signal [990]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[990]) );
  d_ff \sig_prgm_register/genblk1[989].single_DFF  ( .d(
        \sig_prgm_register/or_signal [989]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[989]) );
  d_ff \sig_prgm_register/genblk1[988].single_DFF  ( .d(
        \sig_prgm_register/or_signal [988]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[988]) );
  d_ff \sig_prgm_register/genblk1[987].single_DFF  ( .d(
        \sig_prgm_register/or_signal [987]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[987]) );
  d_ff \sig_prgm_register/genblk1[986].single_DFF  ( .d(
        \sig_prgm_register/or_signal [986]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[986]) );
  d_ff \sig_prgm_register/genblk1[985].single_DFF  ( .d(
        \sig_prgm_register/or_signal [985]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[985]) );
  d_ff \sig_prgm_register/genblk1[984].single_DFF  ( .d(
        \sig_prgm_register/or_signal [984]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[984]) );
  d_ff \sig_prgm_register/genblk1[983].single_DFF  ( .d(
        \sig_prgm_register/or_signal [983]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[983]) );
  d_ff \sig_prgm_register/genblk1[982].single_DFF  ( .d(
        \sig_prgm_register/or_signal [982]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[982]) );
  d_ff \sig_prgm_register/genblk1[981].single_DFF  ( .d(
        \sig_prgm_register/or_signal [981]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[981]) );
  d_ff \sig_prgm_register/genblk1[980].single_DFF  ( .d(
        \sig_prgm_register/or_signal [980]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[980]) );
  d_ff \sig_prgm_register/genblk1[979].single_DFF  ( .d(
        \sig_prgm_register/or_signal [979]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[979]) );
  d_ff \sig_prgm_register/genblk1[978].single_DFF  ( .d(
        \sig_prgm_register/or_signal [978]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[978]) );
  d_ff \sig_prgm_register/genblk1[977].single_DFF  ( .d(
        \sig_prgm_register/or_signal [977]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[977]) );
  d_ff \sig_prgm_register/genblk1[976].single_DFF  ( .d(
        \sig_prgm_register/or_signal [976]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[976]) );
  d_ff \sig_prgm_register/genblk1[975].single_DFF  ( .d(
        \sig_prgm_register/or_signal [975]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[975]) );
  d_ff \sig_prgm_register/genblk1[974].single_DFF  ( .d(
        \sig_prgm_register/or_signal [974]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[974]) );
  d_ff \sig_prgm_register/genblk1[973].single_DFF  ( .d(
        \sig_prgm_register/or_signal [973]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[973]) );
  d_ff \sig_prgm_register/genblk1[972].single_DFF  ( .d(
        \sig_prgm_register/or_signal [972]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[972]) );
  d_ff \sig_prgm_register/genblk1[971].single_DFF  ( .d(
        \sig_prgm_register/or_signal [971]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[971]) );
  d_ff \sig_prgm_register/genblk1[970].single_DFF  ( .d(
        \sig_prgm_register/or_signal [970]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[970]) );
  d_ff \sig_prgm_register/genblk1[969].single_DFF  ( .d(
        \sig_prgm_register/or_signal [969]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[969]) );
  d_ff \sig_prgm_register/genblk1[968].single_DFF  ( .d(
        \sig_prgm_register/or_signal [968]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[968]) );
  d_ff \sig_prgm_register/genblk1[967].single_DFF  ( .d(
        \sig_prgm_register/or_signal [967]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[967]) );
  d_ff \sig_prgm_register/genblk1[966].single_DFF  ( .d(
        \sig_prgm_register/or_signal [966]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[966]) );
  d_ff \sig_prgm_register/genblk1[965].single_DFF  ( .d(
        \sig_prgm_register/or_signal [965]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[965]) );
  d_ff \sig_prgm_register/genblk1[964].single_DFF  ( .d(
        \sig_prgm_register/or_signal [964]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[964]) );
  d_ff \sig_prgm_register/genblk1[963].single_DFF  ( .d(
        \sig_prgm_register/or_signal [963]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[963]) );
  d_ff \sig_prgm_register/genblk1[962].single_DFF  ( .d(
        \sig_prgm_register/or_signal [962]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[962]) );
  d_ff \sig_prgm_register/genblk1[961].single_DFF  ( .d(
        \sig_prgm_register/or_signal [961]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[961]) );
  d_ff \sig_prgm_register/genblk1[960].single_DFF  ( .d(
        \sig_prgm_register/or_signal [960]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[960]) );
  d_ff \sig_prgm_register/genblk1[959].single_DFF  ( .d(
        \sig_prgm_register/or_signal [959]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[959]) );
  d_ff \sig_prgm_register/genblk1[958].single_DFF  ( .d(
        \sig_prgm_register/or_signal [958]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[958]) );
  d_ff \sig_prgm_register/genblk1[957].single_DFF  ( .d(
        \sig_prgm_register/or_signal [957]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[957]) );
  d_ff \sig_prgm_register/genblk1[956].single_DFF  ( .d(
        \sig_prgm_register/or_signal [956]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[956]) );
  d_ff \sig_prgm_register/genblk1[955].single_DFF  ( .d(
        \sig_prgm_register/or_signal [955]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[955]) );
  d_ff \sig_prgm_register/genblk1[954].single_DFF  ( .d(
        \sig_prgm_register/or_signal [954]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[954]) );
  d_ff \sig_prgm_register/genblk1[953].single_DFF  ( .d(
        \sig_prgm_register/or_signal [953]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[953]) );
  d_ff \sig_prgm_register/genblk1[952].single_DFF  ( .d(
        \sig_prgm_register/or_signal [952]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[952]) );
  d_ff \sig_prgm_register/genblk1[951].single_DFF  ( .d(
        \sig_prgm_register/or_signal [951]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[951]) );
  d_ff \sig_prgm_register/genblk1[950].single_DFF  ( .d(
        \sig_prgm_register/or_signal [950]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[950]) );
  d_ff \sig_prgm_register/genblk1[949].single_DFF  ( .d(
        \sig_prgm_register/or_signal [949]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[949]) );
  d_ff \sig_prgm_register/genblk1[948].single_DFF  ( .d(
        \sig_prgm_register/or_signal [948]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[948]) );
  d_ff \sig_prgm_register/genblk1[947].single_DFF  ( .d(
        \sig_prgm_register/or_signal [947]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[947]) );
  d_ff \sig_prgm_register/genblk1[946].single_DFF  ( .d(
        \sig_prgm_register/or_signal [946]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[946]) );
  d_ff \sig_prgm_register/genblk1[945].single_DFF  ( .d(
        \sig_prgm_register/or_signal [945]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[945]) );
  d_ff \sig_prgm_register/genblk1[944].single_DFF  ( .d(
        \sig_prgm_register/or_signal [944]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[944]) );
  d_ff \sig_prgm_register/genblk1[943].single_DFF  ( .d(
        \sig_prgm_register/or_signal [943]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[943]) );
  d_ff \sig_prgm_register/genblk1[942].single_DFF  ( .d(
        \sig_prgm_register/or_signal [942]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[942]) );
  d_ff \sig_prgm_register/genblk1[941].single_DFF  ( .d(
        \sig_prgm_register/or_signal [941]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[941]) );
  d_ff \sig_prgm_register/genblk1[940].single_DFF  ( .d(
        \sig_prgm_register/or_signal [940]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[940]) );
  d_ff \sig_prgm_register/genblk1[939].single_DFF  ( .d(
        \sig_prgm_register/or_signal [939]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[939]) );
  d_ff \sig_prgm_register/genblk1[938].single_DFF  ( .d(
        \sig_prgm_register/or_signal [938]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[938]) );
  d_ff \sig_prgm_register/genblk1[937].single_DFF  ( .d(
        \sig_prgm_register/or_signal [937]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[937]) );
  d_ff \sig_prgm_register/genblk1[936].single_DFF  ( .d(
        \sig_prgm_register/or_signal [936]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[936]) );
  d_ff \sig_prgm_register/genblk1[935].single_DFF  ( .d(
        \sig_prgm_register/or_signal [935]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[935]) );
  d_ff \sig_prgm_register/genblk1[934].single_DFF  ( .d(
        \sig_prgm_register/or_signal [934]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[934]) );
  d_ff \sig_prgm_register/genblk1[933].single_DFF  ( .d(
        \sig_prgm_register/or_signal [933]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[933]) );
  d_ff \sig_prgm_register/genblk1[932].single_DFF  ( .d(
        \sig_prgm_register/or_signal [932]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[932]) );
  d_ff \sig_prgm_register/genblk1[931].single_DFF  ( .d(
        \sig_prgm_register/or_signal [931]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[931]) );
  d_ff \sig_prgm_register/genblk1[930].single_DFF  ( .d(
        \sig_prgm_register/or_signal [930]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[930]) );
  d_ff \sig_prgm_register/genblk1[929].single_DFF  ( .d(
        \sig_prgm_register/or_signal [929]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[929]) );
  d_ff \sig_prgm_register/genblk1[928].single_DFF  ( .d(
        \sig_prgm_register/or_signal [928]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[928]) );
  d_ff \sig_prgm_register/genblk1[927].single_DFF  ( .d(
        \sig_prgm_register/or_signal [927]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[927]) );
  d_ff \sig_prgm_register/genblk1[926].single_DFF  ( .d(
        \sig_prgm_register/or_signal [926]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[926]) );
  d_ff \sig_prgm_register/genblk1[925].single_DFF  ( .d(
        \sig_prgm_register/or_signal [925]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[925]) );
  d_ff \sig_prgm_register/genblk1[924].single_DFF  ( .d(
        \sig_prgm_register/or_signal [924]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[924]) );
  d_ff \sig_prgm_register/genblk1[923].single_DFF  ( .d(
        \sig_prgm_register/or_signal [923]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[923]) );
  d_ff \sig_prgm_register/genblk1[922].single_DFF  ( .d(
        \sig_prgm_register/or_signal [922]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[922]) );
  d_ff \sig_prgm_register/genblk1[921].single_DFF  ( .d(
        \sig_prgm_register/or_signal [921]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[921]) );
  d_ff \sig_prgm_register/genblk1[920].single_DFF  ( .d(
        \sig_prgm_register/or_signal [920]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[920]) );
  d_ff \sig_prgm_register/genblk1[919].single_DFF  ( .d(
        \sig_prgm_register/or_signal [919]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[919]) );
  d_ff \sig_prgm_register/genblk1[918].single_DFF  ( .d(
        \sig_prgm_register/or_signal [918]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[918]) );
  d_ff \sig_prgm_register/genblk1[917].single_DFF  ( .d(
        \sig_prgm_register/or_signal [917]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[917]) );
  d_ff \sig_prgm_register/genblk1[916].single_DFF  ( .d(
        \sig_prgm_register/or_signal [916]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[916]) );
  d_ff \sig_prgm_register/genblk1[915].single_DFF  ( .d(
        \sig_prgm_register/or_signal [915]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[915]) );
  d_ff \sig_prgm_register/genblk1[914].single_DFF  ( .d(
        \sig_prgm_register/or_signal [914]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[914]) );
  d_ff \sig_prgm_register/genblk1[913].single_DFF  ( .d(
        \sig_prgm_register/or_signal [913]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[913]) );
  d_ff \sig_prgm_register/genblk1[912].single_DFF  ( .d(
        \sig_prgm_register/or_signal [912]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[912]) );
  d_ff \sig_prgm_register/genblk1[911].single_DFF  ( .d(
        \sig_prgm_register/or_signal [911]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[911]) );
  d_ff \sig_prgm_register/genblk1[910].single_DFF  ( .d(
        \sig_prgm_register/or_signal [910]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[910]) );
  d_ff \sig_prgm_register/genblk1[909].single_DFF  ( .d(
        \sig_prgm_register/or_signal [909]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[909]) );
  d_ff \sig_prgm_register/genblk1[908].single_DFF  ( .d(
        \sig_prgm_register/or_signal [908]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[908]) );
  d_ff \sig_prgm_register/genblk1[907].single_DFF  ( .d(
        \sig_prgm_register/or_signal [907]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[907]) );
  d_ff \sig_prgm_register/genblk1[906].single_DFF  ( .d(
        \sig_prgm_register/or_signal [906]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[906]) );
  d_ff \sig_prgm_register/genblk1[905].single_DFF  ( .d(
        \sig_prgm_register/or_signal [905]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[905]) );
  d_ff \sig_prgm_register/genblk1[904].single_DFF  ( .d(
        \sig_prgm_register/or_signal [904]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[904]) );
  d_ff \sig_prgm_register/genblk1[903].single_DFF  ( .d(
        \sig_prgm_register/or_signal [903]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[903]) );
  d_ff \sig_prgm_register/genblk1[902].single_DFF  ( .d(
        \sig_prgm_register/or_signal [902]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[902]) );
  d_ff \sig_prgm_register/genblk1[901].single_DFF  ( .d(
        \sig_prgm_register/or_signal [901]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[901]) );
  d_ff \sig_prgm_register/genblk1[900].single_DFF  ( .d(
        \sig_prgm_register/or_signal [900]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[900]) );
  d_ff \sig_prgm_register/genblk1[899].single_DFF  ( .d(
        \sig_prgm_register/or_signal [899]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[899]) );
  d_ff \sig_prgm_register/genblk1[898].single_DFF  ( .d(
        \sig_prgm_register/or_signal [898]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[898]) );
  d_ff \sig_prgm_register/genblk1[897].single_DFF  ( .d(
        \sig_prgm_register/or_signal [897]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[897]) );
  d_ff \sig_prgm_register/genblk1[896].single_DFF  ( .d(
        \sig_prgm_register/or_signal [896]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[896]) );
  d_ff \sig_prgm_register/genblk1[895].single_DFF  ( .d(
        \sig_prgm_register/or_signal [895]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[895]) );
  d_ff \sig_prgm_register/genblk1[894].single_DFF  ( .d(
        \sig_prgm_register/or_signal [894]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[894]) );
  d_ff \sig_prgm_register/genblk1[893].single_DFF  ( .d(
        \sig_prgm_register/or_signal [893]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[893]) );
  d_ff \sig_prgm_register/genblk1[892].single_DFF  ( .d(
        \sig_prgm_register/or_signal [892]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[892]) );
  d_ff \sig_prgm_register/genblk1[891].single_DFF  ( .d(
        \sig_prgm_register/or_signal [891]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[891]) );
  d_ff \sig_prgm_register/genblk1[890].single_DFF  ( .d(
        \sig_prgm_register/or_signal [890]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[890]) );
  d_ff \sig_prgm_register/genblk1[889].single_DFF  ( .d(
        \sig_prgm_register/or_signal [889]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[889]) );
  d_ff \sig_prgm_register/genblk1[888].single_DFF  ( .d(
        \sig_prgm_register/or_signal [888]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[888]) );
  d_ff \sig_prgm_register/genblk1[887].single_DFF  ( .d(
        \sig_prgm_register/or_signal [887]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[887]) );
  d_ff \sig_prgm_register/genblk1[886].single_DFF  ( .d(
        \sig_prgm_register/or_signal [886]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[886]) );
  d_ff \sig_prgm_register/genblk1[885].single_DFF  ( .d(
        \sig_prgm_register/or_signal [885]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[885]) );
  d_ff \sig_prgm_register/genblk1[884].single_DFF  ( .d(
        \sig_prgm_register/or_signal [884]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[884]) );
  d_ff \sig_prgm_register/genblk1[883].single_DFF  ( .d(
        \sig_prgm_register/or_signal [883]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[883]) );
  d_ff \sig_prgm_register/genblk1[882].single_DFF  ( .d(
        \sig_prgm_register/or_signal [882]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[882]) );
  d_ff \sig_prgm_register/genblk1[881].single_DFF  ( .d(
        \sig_prgm_register/or_signal [881]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[881]) );
  d_ff \sig_prgm_register/genblk1[880].single_DFF  ( .d(
        \sig_prgm_register/or_signal [880]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[880]) );
  d_ff \sig_prgm_register/genblk1[879].single_DFF  ( .d(
        \sig_prgm_register/or_signal [879]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[879]) );
  d_ff \sig_prgm_register/genblk1[878].single_DFF  ( .d(
        \sig_prgm_register/or_signal [878]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[878]) );
  d_ff \sig_prgm_register/genblk1[877].single_DFF  ( .d(
        \sig_prgm_register/or_signal [877]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[877]) );
  d_ff \sig_prgm_register/genblk1[876].single_DFF  ( .d(
        \sig_prgm_register/or_signal [876]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[876]) );
  d_ff \sig_prgm_register/genblk1[875].single_DFF  ( .d(
        \sig_prgm_register/or_signal [875]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[875]) );
  d_ff \sig_prgm_register/genblk1[874].single_DFF  ( .d(
        \sig_prgm_register/or_signal [874]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[874]) );
  d_ff \sig_prgm_register/genblk1[873].single_DFF  ( .d(
        \sig_prgm_register/or_signal [873]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[873]) );
  d_ff \sig_prgm_register/genblk1[872].single_DFF  ( .d(
        \sig_prgm_register/or_signal [872]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[872]) );
  d_ff \sig_prgm_register/genblk1[871].single_DFF  ( .d(
        \sig_prgm_register/or_signal [871]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[871]) );
  d_ff \sig_prgm_register/genblk1[870].single_DFF  ( .d(
        \sig_prgm_register/or_signal [870]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[870]) );
  d_ff \sig_prgm_register/genblk1[869].single_DFF  ( .d(
        \sig_prgm_register/or_signal [869]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[869]) );
  d_ff \sig_prgm_register/genblk1[868].single_DFF  ( .d(
        \sig_prgm_register/or_signal [868]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[868]) );
  d_ff \sig_prgm_register/genblk1[867].single_DFF  ( .d(
        \sig_prgm_register/or_signal [867]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[867]) );
  d_ff \sig_prgm_register/genblk1[866].single_DFF  ( .d(
        \sig_prgm_register/or_signal [866]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[866]) );
  d_ff \sig_prgm_register/genblk1[865].single_DFF  ( .d(
        \sig_prgm_register/or_signal [865]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[865]) );
  d_ff \sig_prgm_register/genblk1[864].single_DFF  ( .d(
        \sig_prgm_register/or_signal [864]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[864]) );
  d_ff \sig_prgm_register/genblk1[863].single_DFF  ( .d(
        \sig_prgm_register/or_signal [863]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[863]) );
  d_ff \sig_prgm_register/genblk1[862].single_DFF  ( .d(
        \sig_prgm_register/or_signal [862]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[862]) );
  d_ff \sig_prgm_register/genblk1[861].single_DFF  ( .d(
        \sig_prgm_register/or_signal [861]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[861]) );
  d_ff \sig_prgm_register/genblk1[860].single_DFF  ( .d(
        \sig_prgm_register/or_signal [860]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[860]) );
  d_ff \sig_prgm_register/genblk1[859].single_DFF  ( .d(
        \sig_prgm_register/or_signal [859]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[859]) );
  d_ff \sig_prgm_register/genblk1[858].single_DFF  ( .d(
        \sig_prgm_register/or_signal [858]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[858]) );
  d_ff \sig_prgm_register/genblk1[857].single_DFF  ( .d(
        \sig_prgm_register/or_signal [857]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[857]) );
  d_ff \sig_prgm_register/genblk1[856].single_DFF  ( .d(
        \sig_prgm_register/or_signal [856]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[856]) );
  d_ff \sig_prgm_register/genblk1[855].single_DFF  ( .d(
        \sig_prgm_register/or_signal [855]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[855]) );
  d_ff \sig_prgm_register/genblk1[854].single_DFF  ( .d(
        \sig_prgm_register/or_signal [854]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[854]) );
  d_ff \sig_prgm_register/genblk1[853].single_DFF  ( .d(
        \sig_prgm_register/or_signal [853]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[853]) );
  d_ff \sig_prgm_register/genblk1[852].single_DFF  ( .d(
        \sig_prgm_register/or_signal [852]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[852]) );
  d_ff \sig_prgm_register/genblk1[851].single_DFF  ( .d(
        \sig_prgm_register/or_signal [851]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[851]) );
  d_ff \sig_prgm_register/genblk1[850].single_DFF  ( .d(
        \sig_prgm_register/or_signal [850]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[850]) );
  d_ff \sig_prgm_register/genblk1[849].single_DFF  ( .d(
        \sig_prgm_register/or_signal [849]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[849]) );
  d_ff \sig_prgm_register/genblk1[848].single_DFF  ( .d(
        \sig_prgm_register/or_signal [848]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[848]) );
  d_ff \sig_prgm_register/genblk1[847].single_DFF  ( .d(
        \sig_prgm_register/or_signal [847]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[847]) );
  d_ff \sig_prgm_register/genblk1[846].single_DFF  ( .d(
        \sig_prgm_register/or_signal [846]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[846]) );
  d_ff \sig_prgm_register/genblk1[845].single_DFF  ( .d(
        \sig_prgm_register/or_signal [845]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[845]) );
  d_ff \sig_prgm_register/genblk1[844].single_DFF  ( .d(
        \sig_prgm_register/or_signal [844]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[844]) );
  d_ff \sig_prgm_register/genblk1[843].single_DFF  ( .d(
        \sig_prgm_register/or_signal [843]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[843]) );
  d_ff \sig_prgm_register/genblk1[842].single_DFF  ( .d(
        \sig_prgm_register/or_signal [842]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[842]) );
  d_ff \sig_prgm_register/genblk1[841].single_DFF  ( .d(
        \sig_prgm_register/or_signal [841]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[841]) );
  d_ff \sig_prgm_register/genblk1[840].single_DFF  ( .d(
        \sig_prgm_register/or_signal [840]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[840]) );
  d_ff \sig_prgm_register/genblk1[839].single_DFF  ( .d(
        \sig_prgm_register/or_signal [839]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[839]) );
  d_ff \sig_prgm_register/genblk1[838].single_DFF  ( .d(
        \sig_prgm_register/or_signal [838]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[838]) );
  d_ff \sig_prgm_register/genblk1[837].single_DFF  ( .d(
        \sig_prgm_register/or_signal [837]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[837]) );
  d_ff \sig_prgm_register/genblk1[836].single_DFF  ( .d(
        \sig_prgm_register/or_signal [836]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[836]) );
  d_ff \sig_prgm_register/genblk1[835].single_DFF  ( .d(
        \sig_prgm_register/or_signal [835]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[835]) );
  d_ff \sig_prgm_register/genblk1[834].single_DFF  ( .d(
        \sig_prgm_register/or_signal [834]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[834]) );
  d_ff \sig_prgm_register/genblk1[833].single_DFF  ( .d(
        \sig_prgm_register/or_signal [833]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[833]) );
  d_ff \sig_prgm_register/genblk1[832].single_DFF  ( .d(
        \sig_prgm_register/or_signal [832]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[832]) );
  d_ff \sig_prgm_register/genblk1[831].single_DFF  ( .d(
        \sig_prgm_register/or_signal [831]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[831]) );
  d_ff \sig_prgm_register/genblk1[830].single_DFF  ( .d(
        \sig_prgm_register/or_signal [830]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[830]) );
  d_ff \sig_prgm_register/genblk1[829].single_DFF  ( .d(
        \sig_prgm_register/or_signal [829]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[829]) );
  d_ff \sig_prgm_register/genblk1[828].single_DFF  ( .d(
        \sig_prgm_register/or_signal [828]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[828]) );
  d_ff \sig_prgm_register/genblk1[827].single_DFF  ( .d(
        \sig_prgm_register/or_signal [827]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[827]) );
  d_ff \sig_prgm_register/genblk1[826].single_DFF  ( .d(
        \sig_prgm_register/or_signal [826]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[826]) );
  d_ff \sig_prgm_register/genblk1[825].single_DFF  ( .d(
        \sig_prgm_register/or_signal [825]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[825]) );
  d_ff \sig_prgm_register/genblk1[824].single_DFF  ( .d(
        \sig_prgm_register/or_signal [824]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[824]) );
  d_ff \sig_prgm_register/genblk1[823].single_DFF  ( .d(
        \sig_prgm_register/or_signal [823]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[823]) );
  d_ff \sig_prgm_register/genblk1[822].single_DFF  ( .d(
        \sig_prgm_register/or_signal [822]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[822]) );
  d_ff \sig_prgm_register/genblk1[821].single_DFF  ( .d(
        \sig_prgm_register/or_signal [821]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[821]) );
  d_ff \sig_prgm_register/genblk1[820].single_DFF  ( .d(
        \sig_prgm_register/or_signal [820]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[820]) );
  d_ff \sig_prgm_register/genblk1[819].single_DFF  ( .d(
        \sig_prgm_register/or_signal [819]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[819]) );
  d_ff \sig_prgm_register/genblk1[818].single_DFF  ( .d(
        \sig_prgm_register/or_signal [818]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[818]) );
  d_ff \sig_prgm_register/genblk1[817].single_DFF  ( .d(
        \sig_prgm_register/or_signal [817]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[817]) );
  d_ff \sig_prgm_register/genblk1[816].single_DFF  ( .d(
        \sig_prgm_register/or_signal [816]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[816]) );
  d_ff \sig_prgm_register/genblk1[815].single_DFF  ( .d(
        \sig_prgm_register/or_signal [815]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[815]) );
  d_ff \sig_prgm_register/genblk1[814].single_DFF  ( .d(
        \sig_prgm_register/or_signal [814]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[814]) );
  d_ff \sig_prgm_register/genblk1[813].single_DFF  ( .d(
        \sig_prgm_register/or_signal [813]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[813]) );
  d_ff \sig_prgm_register/genblk1[812].single_DFF  ( .d(
        \sig_prgm_register/or_signal [812]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[812]) );
  d_ff \sig_prgm_register/genblk1[811].single_DFF  ( .d(
        \sig_prgm_register/or_signal [811]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[811]) );
  d_ff \sig_prgm_register/genblk1[810].single_DFF  ( .d(
        \sig_prgm_register/or_signal [810]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[810]) );
  d_ff \sig_prgm_register/genblk1[809].single_DFF  ( .d(
        \sig_prgm_register/or_signal [809]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[809]) );
  d_ff \sig_prgm_register/genblk1[808].single_DFF  ( .d(
        \sig_prgm_register/or_signal [808]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[808]) );
  d_ff \sig_prgm_register/genblk1[807].single_DFF  ( .d(
        \sig_prgm_register/or_signal [807]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[807]) );
  d_ff \sig_prgm_register/genblk1[806].single_DFF  ( .d(
        \sig_prgm_register/or_signal [806]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[806]) );
  d_ff \sig_prgm_register/genblk1[805].single_DFF  ( .d(
        \sig_prgm_register/or_signal [805]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[805]) );
  d_ff \sig_prgm_register/genblk1[804].single_DFF  ( .d(
        \sig_prgm_register/or_signal [804]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[804]) );
  d_ff \sig_prgm_register/genblk1[803].single_DFF  ( .d(
        \sig_prgm_register/or_signal [803]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[803]) );
  d_ff \sig_prgm_register/genblk1[802].single_DFF  ( .d(
        \sig_prgm_register/or_signal [802]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[802]) );
  d_ff \sig_prgm_register/genblk1[801].single_DFF  ( .d(
        \sig_prgm_register/or_signal [801]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[801]) );
  d_ff \sig_prgm_register/genblk1[800].single_DFF  ( .d(
        \sig_prgm_register/or_signal [800]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[800]) );
  d_ff \sig_prgm_register/genblk1[799].single_DFF  ( .d(
        \sig_prgm_register/or_signal [799]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[799]) );
  d_ff \sig_prgm_register/genblk1[798].single_DFF  ( .d(
        \sig_prgm_register/or_signal [798]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[798]) );
  d_ff \sig_prgm_register/genblk1[797].single_DFF  ( .d(
        \sig_prgm_register/or_signal [797]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[797]) );
  d_ff \sig_prgm_register/genblk1[796].single_DFF  ( .d(
        \sig_prgm_register/or_signal [796]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[796]) );
  d_ff \sig_prgm_register/genblk1[795].single_DFF  ( .d(
        \sig_prgm_register/or_signal [795]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[795]) );
  d_ff \sig_prgm_register/genblk1[794].single_DFF  ( .d(
        \sig_prgm_register/or_signal [794]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[794]) );
  d_ff \sig_prgm_register/genblk1[793].single_DFF  ( .d(
        \sig_prgm_register/or_signal [793]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[793]) );
  d_ff \sig_prgm_register/genblk1[792].single_DFF  ( .d(
        \sig_prgm_register/or_signal [792]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[792]) );
  d_ff \sig_prgm_register/genblk1[791].single_DFF  ( .d(
        \sig_prgm_register/or_signal [791]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[791]) );
  d_ff \sig_prgm_register/genblk1[790].single_DFF  ( .d(
        \sig_prgm_register/or_signal [790]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[790]) );
  d_ff \sig_prgm_register/genblk1[789].single_DFF  ( .d(
        \sig_prgm_register/or_signal [789]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[789]) );
  d_ff \sig_prgm_register/genblk1[788].single_DFF  ( .d(
        \sig_prgm_register/or_signal [788]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[788]) );
  d_ff \sig_prgm_register/genblk1[787].single_DFF  ( .d(
        \sig_prgm_register/or_signal [787]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[787]) );
  d_ff \sig_prgm_register/genblk1[786].single_DFF  ( .d(
        \sig_prgm_register/or_signal [786]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[786]) );
  d_ff \sig_prgm_register/genblk1[785].single_DFF  ( .d(
        \sig_prgm_register/or_signal [785]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[785]) );
  d_ff \sig_prgm_register/genblk1[784].single_DFF  ( .d(
        \sig_prgm_register/or_signal [784]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[784]) );
  d_ff \sig_prgm_register/genblk1[783].single_DFF  ( .d(
        \sig_prgm_register/or_signal [783]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[783]) );
  d_ff \sig_prgm_register/genblk1[782].single_DFF  ( .d(
        \sig_prgm_register/or_signal [782]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[782]) );
  d_ff \sig_prgm_register/genblk1[781].single_DFF  ( .d(
        \sig_prgm_register/or_signal [781]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[781]) );
  d_ff \sig_prgm_register/genblk1[780].single_DFF  ( .d(
        \sig_prgm_register/or_signal [780]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[780]) );
  d_ff \sig_prgm_register/genblk1[779].single_DFF  ( .d(
        \sig_prgm_register/or_signal [779]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[779]) );
  d_ff \sig_prgm_register/genblk1[778].single_DFF  ( .d(
        \sig_prgm_register/or_signal [778]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[778]) );
  d_ff \sig_prgm_register/genblk1[777].single_DFF  ( .d(
        \sig_prgm_register/or_signal [777]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[777]) );
  d_ff \sig_prgm_register/genblk1[776].single_DFF  ( .d(
        \sig_prgm_register/or_signal [776]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[776]) );
  d_ff \sig_prgm_register/genblk1[775].single_DFF  ( .d(
        \sig_prgm_register/or_signal [775]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[775]) );
  d_ff \sig_prgm_register/genblk1[774].single_DFF  ( .d(
        \sig_prgm_register/or_signal [774]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[774]) );
  d_ff \sig_prgm_register/genblk1[773].single_DFF  ( .d(
        \sig_prgm_register/or_signal [773]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[773]) );
  d_ff \sig_prgm_register/genblk1[772].single_DFF  ( .d(
        \sig_prgm_register/or_signal [772]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[772]) );
  d_ff \sig_prgm_register/genblk1[771].single_DFF  ( .d(
        \sig_prgm_register/or_signal [771]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[771]) );
  d_ff \sig_prgm_register/genblk1[770].single_DFF  ( .d(
        \sig_prgm_register/or_signal [770]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[770]) );
  d_ff \sig_prgm_register/genblk1[769].single_DFF  ( .d(
        \sig_prgm_register/or_signal [769]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[769]) );
  d_ff \sig_prgm_register/genblk1[768].single_DFF  ( .d(
        \sig_prgm_register/or_signal [768]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[768]) );
  d_ff \sig_prgm_register/genblk1[767].single_DFF  ( .d(
        \sig_prgm_register/or_signal [767]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[767]) );
  d_ff \sig_prgm_register/genblk1[766].single_DFF  ( .d(
        \sig_prgm_register/or_signal [766]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[766]) );
  d_ff \sig_prgm_register/genblk1[765].single_DFF  ( .d(
        \sig_prgm_register/or_signal [765]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[765]) );
  d_ff \sig_prgm_register/genblk1[764].single_DFF  ( .d(
        \sig_prgm_register/or_signal [764]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[764]) );
  d_ff \sig_prgm_register/genblk1[763].single_DFF  ( .d(
        \sig_prgm_register/or_signal [763]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[763]) );
  d_ff \sig_prgm_register/genblk1[762].single_DFF  ( .d(
        \sig_prgm_register/or_signal [762]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[762]) );
  d_ff \sig_prgm_register/genblk1[761].single_DFF  ( .d(
        \sig_prgm_register/or_signal [761]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[761]) );
  d_ff \sig_prgm_register/genblk1[760].single_DFF  ( .d(
        \sig_prgm_register/or_signal [760]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[760]) );
  d_ff \sig_prgm_register/genblk1[759].single_DFF  ( .d(
        \sig_prgm_register/or_signal [759]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[759]) );
  d_ff \sig_prgm_register/genblk1[758].single_DFF  ( .d(
        \sig_prgm_register/or_signal [758]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[758]) );
  d_ff \sig_prgm_register/genblk1[757].single_DFF  ( .d(
        \sig_prgm_register/or_signal [757]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[757]) );
  d_ff \sig_prgm_register/genblk1[756].single_DFF  ( .d(
        \sig_prgm_register/or_signal [756]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[756]) );
  d_ff \sig_prgm_register/genblk1[755].single_DFF  ( .d(
        \sig_prgm_register/or_signal [755]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[755]) );
  d_ff \sig_prgm_register/genblk1[754].single_DFF  ( .d(
        \sig_prgm_register/or_signal [754]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[754]) );
  d_ff \sig_prgm_register/genblk1[753].single_DFF  ( .d(
        \sig_prgm_register/or_signal [753]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[753]) );
  d_ff \sig_prgm_register/genblk1[752].single_DFF  ( .d(
        \sig_prgm_register/or_signal [752]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[752]) );
  d_ff \sig_prgm_register/genblk1[751].single_DFF  ( .d(
        \sig_prgm_register/or_signal [751]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[751]) );
  d_ff \sig_prgm_register/genblk1[750].single_DFF  ( .d(
        \sig_prgm_register/or_signal [750]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[750]) );
  d_ff \sig_prgm_register/genblk1[749].single_DFF  ( .d(
        \sig_prgm_register/or_signal [749]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[749]) );
  d_ff \sig_prgm_register/genblk1[748].single_DFF  ( .d(
        \sig_prgm_register/or_signal [748]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[748]) );
  d_ff \sig_prgm_register/genblk1[747].single_DFF  ( .d(
        \sig_prgm_register/or_signal [747]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[747]) );
  d_ff \sig_prgm_register/genblk1[746].single_DFF  ( .d(
        \sig_prgm_register/or_signal [746]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[746]) );
  d_ff \sig_prgm_register/genblk1[745].single_DFF  ( .d(
        \sig_prgm_register/or_signal [745]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[745]) );
  d_ff \sig_prgm_register/genblk1[744].single_DFF  ( .d(
        \sig_prgm_register/or_signal [744]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[744]) );
  d_ff \sig_prgm_register/genblk1[743].single_DFF  ( .d(
        \sig_prgm_register/or_signal [743]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[743]) );
  d_ff \sig_prgm_register/genblk1[742].single_DFF  ( .d(
        \sig_prgm_register/or_signal [742]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[742]) );
  d_ff \sig_prgm_register/genblk1[741].single_DFF  ( .d(
        \sig_prgm_register/or_signal [741]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[741]) );
  d_ff \sig_prgm_register/genblk1[740].single_DFF  ( .d(
        \sig_prgm_register/or_signal [740]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[740]) );
  d_ff \sig_prgm_register/genblk1[739].single_DFF  ( .d(
        \sig_prgm_register/or_signal [739]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[739]) );
  d_ff \sig_prgm_register/genblk1[738].single_DFF  ( .d(
        \sig_prgm_register/or_signal [738]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[738]) );
  d_ff \sig_prgm_register/genblk1[737].single_DFF  ( .d(
        \sig_prgm_register/or_signal [737]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[737]) );
  d_ff \sig_prgm_register/genblk1[736].single_DFF  ( .d(
        \sig_prgm_register/or_signal [736]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[736]) );
  d_ff \sig_prgm_register/genblk1[735].single_DFF  ( .d(
        \sig_prgm_register/or_signal [735]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[735]) );
  d_ff \sig_prgm_register/genblk1[734].single_DFF  ( .d(
        \sig_prgm_register/or_signal [734]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[734]) );
  d_ff \sig_prgm_register/genblk1[733].single_DFF  ( .d(
        \sig_prgm_register/or_signal [733]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[733]) );
  d_ff \sig_prgm_register/genblk1[732].single_DFF  ( .d(
        \sig_prgm_register/or_signal [732]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[732]) );
  d_ff \sig_prgm_register/genblk1[731].single_DFF  ( .d(
        \sig_prgm_register/or_signal [731]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[731]) );
  d_ff \sig_prgm_register/genblk1[730].single_DFF  ( .d(
        \sig_prgm_register/or_signal [730]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[730]) );
  d_ff \sig_prgm_register/genblk1[729].single_DFF  ( .d(
        \sig_prgm_register/or_signal [729]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[729]) );
  d_ff \sig_prgm_register/genblk1[728].single_DFF  ( .d(
        \sig_prgm_register/or_signal [728]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[728]) );
  d_ff \sig_prgm_register/genblk1[727].single_DFF  ( .d(
        \sig_prgm_register/or_signal [727]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[727]) );
  d_ff \sig_prgm_register/genblk1[726].single_DFF  ( .d(
        \sig_prgm_register/or_signal [726]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[726]) );
  d_ff \sig_prgm_register/genblk1[725].single_DFF  ( .d(
        \sig_prgm_register/or_signal [725]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[725]) );
  d_ff \sig_prgm_register/genblk1[724].single_DFF  ( .d(
        \sig_prgm_register/or_signal [724]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[724]) );
  d_ff \sig_prgm_register/genblk1[723].single_DFF  ( .d(
        \sig_prgm_register/or_signal [723]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[723]) );
  d_ff \sig_prgm_register/genblk1[722].single_DFF  ( .d(
        \sig_prgm_register/or_signal [722]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[722]) );
  d_ff \sig_prgm_register/genblk1[721].single_DFF  ( .d(
        \sig_prgm_register/or_signal [721]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[721]) );
  d_ff \sig_prgm_register/genblk1[720].single_DFF  ( .d(
        \sig_prgm_register/or_signal [720]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[720]) );
  d_ff \sig_prgm_register/genblk1[719].single_DFF  ( .d(
        \sig_prgm_register/or_signal [719]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[719]) );
  d_ff \sig_prgm_register/genblk1[718].single_DFF  ( .d(
        \sig_prgm_register/or_signal [718]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[718]) );
  d_ff \sig_prgm_register/genblk1[717].single_DFF  ( .d(
        \sig_prgm_register/or_signal [717]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[717]) );
  d_ff \sig_prgm_register/genblk1[716].single_DFF  ( .d(
        \sig_prgm_register/or_signal [716]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[716]) );
  d_ff \sig_prgm_register/genblk1[715].single_DFF  ( .d(
        \sig_prgm_register/or_signal [715]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[715]) );
  d_ff \sig_prgm_register/genblk1[714].single_DFF  ( .d(
        \sig_prgm_register/or_signal [714]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[714]) );
  d_ff \sig_prgm_register/genblk1[713].single_DFF  ( .d(
        \sig_prgm_register/or_signal [713]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[713]) );
  d_ff \sig_prgm_register/genblk1[712].single_DFF  ( .d(
        \sig_prgm_register/or_signal [712]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[712]) );
  d_ff \sig_prgm_register/genblk1[711].single_DFF  ( .d(
        \sig_prgm_register/or_signal [711]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[711]) );
  d_ff \sig_prgm_register/genblk1[710].single_DFF  ( .d(
        \sig_prgm_register/or_signal [710]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[710]) );
  d_ff \sig_prgm_register/genblk1[709].single_DFF  ( .d(
        \sig_prgm_register/or_signal [709]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[709]) );
  d_ff \sig_prgm_register/genblk1[708].single_DFF  ( .d(
        \sig_prgm_register/or_signal [708]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[708]) );
  d_ff \sig_prgm_register/genblk1[707].single_DFF  ( .d(
        \sig_prgm_register/or_signal [707]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[707]) );
  d_ff \sig_prgm_register/genblk1[706].single_DFF  ( .d(
        \sig_prgm_register/or_signal [706]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[706]) );
  d_ff \sig_prgm_register/genblk1[705].single_DFF  ( .d(
        \sig_prgm_register/or_signal [705]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[705]) );
  d_ff \sig_prgm_register/genblk1[704].single_DFF  ( .d(
        \sig_prgm_register/or_signal [704]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[704]) );
  d_ff \sig_prgm_register/genblk1[703].single_DFF  ( .d(
        \sig_prgm_register/or_signal [703]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[703]) );
  d_ff \sig_prgm_register/genblk1[702].single_DFF  ( .d(
        \sig_prgm_register/or_signal [702]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[702]) );
  d_ff \sig_prgm_register/genblk1[701].single_DFF  ( .d(
        \sig_prgm_register/or_signal [701]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[701]) );
  d_ff \sig_prgm_register/genblk1[700].single_DFF  ( .d(
        \sig_prgm_register/or_signal [700]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[700]) );
  d_ff \sig_prgm_register/genblk1[699].single_DFF  ( .d(
        \sig_prgm_register/or_signal [699]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[699]) );
  d_ff \sig_prgm_register/genblk1[698].single_DFF  ( .d(
        \sig_prgm_register/or_signal [698]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[698]) );
  d_ff \sig_prgm_register/genblk1[697].single_DFF  ( .d(
        \sig_prgm_register/or_signal [697]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[697]) );
  d_ff \sig_prgm_register/genblk1[696].single_DFF  ( .d(
        \sig_prgm_register/or_signal [696]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[696]) );
  d_ff \sig_prgm_register/genblk1[695].single_DFF  ( .d(
        \sig_prgm_register/or_signal [695]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[695]) );
  d_ff \sig_prgm_register/genblk1[694].single_DFF  ( .d(
        \sig_prgm_register/or_signal [694]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[694]) );
  d_ff \sig_prgm_register/genblk1[693].single_DFF  ( .d(
        \sig_prgm_register/or_signal [693]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[693]) );
  d_ff \sig_prgm_register/genblk1[692].single_DFF  ( .d(
        \sig_prgm_register/or_signal [692]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[692]) );
  d_ff \sig_prgm_register/genblk1[691].single_DFF  ( .d(
        \sig_prgm_register/or_signal [691]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[691]) );
  d_ff \sig_prgm_register/genblk1[690].single_DFF  ( .d(
        \sig_prgm_register/or_signal [690]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[690]) );
  d_ff \sig_prgm_register/genblk1[689].single_DFF  ( .d(
        \sig_prgm_register/or_signal [689]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[689]) );
  d_ff \sig_prgm_register/genblk1[688].single_DFF  ( .d(
        \sig_prgm_register/or_signal [688]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[688]) );
  d_ff \sig_prgm_register/genblk1[687].single_DFF  ( .d(
        \sig_prgm_register/or_signal [687]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[687]) );
  d_ff \sig_prgm_register/genblk1[686].single_DFF  ( .d(
        \sig_prgm_register/or_signal [686]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[686]) );
  d_ff \sig_prgm_register/genblk1[685].single_DFF  ( .d(
        \sig_prgm_register/or_signal [685]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[685]) );
  d_ff \sig_prgm_register/genblk1[684].single_DFF  ( .d(
        \sig_prgm_register/or_signal [684]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[684]) );
  d_ff \sig_prgm_register/genblk1[683].single_DFF  ( .d(
        \sig_prgm_register/or_signal [683]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[683]) );
  d_ff \sig_prgm_register/genblk1[682].single_DFF  ( .d(
        \sig_prgm_register/or_signal [682]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[682]) );
  d_ff \sig_prgm_register/genblk1[681].single_DFF  ( .d(
        \sig_prgm_register/or_signal [681]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[681]) );
  d_ff \sig_prgm_register/genblk1[680].single_DFF  ( .d(
        \sig_prgm_register/or_signal [680]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[680]) );
  d_ff \sig_prgm_register/genblk1[679].single_DFF  ( .d(
        \sig_prgm_register/or_signal [679]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[679]) );
  d_ff \sig_prgm_register/genblk1[678].single_DFF  ( .d(
        \sig_prgm_register/or_signal [678]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[678]) );
  d_ff \sig_prgm_register/genblk1[677].single_DFF  ( .d(
        \sig_prgm_register/or_signal [677]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[677]) );
  d_ff \sig_prgm_register/genblk1[676].single_DFF  ( .d(
        \sig_prgm_register/or_signal [676]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[676]) );
  d_ff \sig_prgm_register/genblk1[675].single_DFF  ( .d(
        \sig_prgm_register/or_signal [675]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[675]) );
  d_ff \sig_prgm_register/genblk1[674].single_DFF  ( .d(
        \sig_prgm_register/or_signal [674]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[674]) );
  d_ff \sig_prgm_register/genblk1[673].single_DFF  ( .d(
        \sig_prgm_register/or_signal [673]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[673]) );
  d_ff \sig_prgm_register/genblk1[672].single_DFF  ( .d(
        \sig_prgm_register/or_signal [672]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[672]) );
  d_ff \sig_prgm_register/genblk1[671].single_DFF  ( .d(
        \sig_prgm_register/or_signal [671]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[671]) );
  d_ff \sig_prgm_register/genblk1[670].single_DFF  ( .d(
        \sig_prgm_register/or_signal [670]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[670]) );
  d_ff \sig_prgm_register/genblk1[669].single_DFF  ( .d(
        \sig_prgm_register/or_signal [669]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[669]) );
  d_ff \sig_prgm_register/genblk1[668].single_DFF  ( .d(
        \sig_prgm_register/or_signal [668]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[668]) );
  d_ff \sig_prgm_register/genblk1[667].single_DFF  ( .d(
        \sig_prgm_register/or_signal [667]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[667]) );
  d_ff \sig_prgm_register/genblk1[666].single_DFF  ( .d(
        \sig_prgm_register/or_signal [666]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[666]) );
  d_ff \sig_prgm_register/genblk1[665].single_DFF  ( .d(
        \sig_prgm_register/or_signal [665]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[665]) );
  d_ff \sig_prgm_register/genblk1[664].single_DFF  ( .d(
        \sig_prgm_register/or_signal [664]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[664]) );
  d_ff \sig_prgm_register/genblk1[663].single_DFF  ( .d(
        \sig_prgm_register/or_signal [663]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[663]) );
  d_ff \sig_prgm_register/genblk1[662].single_DFF  ( .d(
        \sig_prgm_register/or_signal [662]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[662]) );
  d_ff \sig_prgm_register/genblk1[661].single_DFF  ( .d(
        \sig_prgm_register/or_signal [661]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[661]) );
  d_ff \sig_prgm_register/genblk1[660].single_DFF  ( .d(
        \sig_prgm_register/or_signal [660]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[660]) );
  d_ff \sig_prgm_register/genblk1[659].single_DFF  ( .d(
        \sig_prgm_register/or_signal [659]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[659]) );
  d_ff \sig_prgm_register/genblk1[658].single_DFF  ( .d(
        \sig_prgm_register/or_signal [658]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[658]) );
  d_ff \sig_prgm_register/genblk1[657].single_DFF  ( .d(
        \sig_prgm_register/or_signal [657]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[657]) );
  d_ff \sig_prgm_register/genblk1[656].single_DFF  ( .d(
        \sig_prgm_register/or_signal [656]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[656]) );
  d_ff \sig_prgm_register/genblk1[655].single_DFF  ( .d(
        \sig_prgm_register/or_signal [655]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[655]) );
  d_ff \sig_prgm_register/genblk1[654].single_DFF  ( .d(
        \sig_prgm_register/or_signal [654]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[654]) );
  d_ff \sig_prgm_register/genblk1[653].single_DFF  ( .d(
        \sig_prgm_register/or_signal [653]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[653]) );
  d_ff \sig_prgm_register/genblk1[652].single_DFF  ( .d(
        \sig_prgm_register/or_signal [652]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[652]) );
  d_ff \sig_prgm_register/genblk1[651].single_DFF  ( .d(
        \sig_prgm_register/or_signal [651]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[651]) );
  d_ff \sig_prgm_register/genblk1[650].single_DFF  ( .d(
        \sig_prgm_register/or_signal [650]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[650]) );
  d_ff \sig_prgm_register/genblk1[649].single_DFF  ( .d(
        \sig_prgm_register/or_signal [649]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[649]) );
  d_ff \sig_prgm_register/genblk1[648].single_DFF  ( .d(
        \sig_prgm_register/or_signal [648]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[648]) );
  d_ff \sig_prgm_register/genblk1[647].single_DFF  ( .d(
        \sig_prgm_register/or_signal [647]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[647]) );
  d_ff \sig_prgm_register/genblk1[646].single_DFF  ( .d(
        \sig_prgm_register/or_signal [646]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[646]) );
  d_ff \sig_prgm_register/genblk1[645].single_DFF  ( .d(
        \sig_prgm_register/or_signal [645]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[645]) );
  d_ff \sig_prgm_register/genblk1[644].single_DFF  ( .d(
        \sig_prgm_register/or_signal [644]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[644]) );
  d_ff \sig_prgm_register/genblk1[643].single_DFF  ( .d(
        \sig_prgm_register/or_signal [643]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[643]) );
  d_ff \sig_prgm_register/genblk1[642].single_DFF  ( .d(
        \sig_prgm_register/or_signal [642]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[642]) );
  d_ff \sig_prgm_register/genblk1[641].single_DFF  ( .d(
        \sig_prgm_register/or_signal [641]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[641]) );
  d_ff \sig_prgm_register/genblk1[640].single_DFF  ( .d(
        \sig_prgm_register/or_signal [640]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[640]) );
  d_ff \sig_prgm_register/genblk1[639].single_DFF  ( .d(
        \sig_prgm_register/or_signal [639]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[639]) );
  d_ff \sig_prgm_register/genblk1[638].single_DFF  ( .d(
        \sig_prgm_register/or_signal [638]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[638]) );
  d_ff \sig_prgm_register/genblk1[637].single_DFF  ( .d(
        \sig_prgm_register/or_signal [637]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[637]) );
  d_ff \sig_prgm_register/genblk1[636].single_DFF  ( .d(
        \sig_prgm_register/or_signal [636]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[636]) );
  d_ff \sig_prgm_register/genblk1[635].single_DFF  ( .d(
        \sig_prgm_register/or_signal [635]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[635]) );
  d_ff \sig_prgm_register/genblk1[634].single_DFF  ( .d(
        \sig_prgm_register/or_signal [634]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[634]) );
  d_ff \sig_prgm_register/genblk1[633].single_DFF  ( .d(
        \sig_prgm_register/or_signal [633]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[633]) );
  d_ff \sig_prgm_register/genblk1[632].single_DFF  ( .d(
        \sig_prgm_register/or_signal [632]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[632]) );
  d_ff \sig_prgm_register/genblk1[631].single_DFF  ( .d(
        \sig_prgm_register/or_signal [631]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[631]) );
  d_ff \sig_prgm_register/genblk1[630].single_DFF  ( .d(
        \sig_prgm_register/or_signal [630]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[630]) );
  d_ff \sig_prgm_register/genblk1[629].single_DFF  ( .d(
        \sig_prgm_register/or_signal [629]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[629]) );
  d_ff \sig_prgm_register/genblk1[628].single_DFF  ( .d(
        \sig_prgm_register/or_signal [628]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[628]) );
  d_ff \sig_prgm_register/genblk1[627].single_DFF  ( .d(
        \sig_prgm_register/or_signal [627]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[627]) );
  d_ff \sig_prgm_register/genblk1[626].single_DFF  ( .d(
        \sig_prgm_register/or_signal [626]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[626]) );
  d_ff \sig_prgm_register/genblk1[625].single_DFF  ( .d(
        \sig_prgm_register/or_signal [625]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[625]) );
  d_ff \sig_prgm_register/genblk1[624].single_DFF  ( .d(
        \sig_prgm_register/or_signal [624]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[624]) );
  d_ff \sig_prgm_register/genblk1[623].single_DFF  ( .d(
        \sig_prgm_register/or_signal [623]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[623]) );
  d_ff \sig_prgm_register/genblk1[622].single_DFF  ( .d(
        \sig_prgm_register/or_signal [622]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[622]) );
  d_ff \sig_prgm_register/genblk1[621].single_DFF  ( .d(
        \sig_prgm_register/or_signal [621]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[621]) );
  d_ff \sig_prgm_register/genblk1[620].single_DFF  ( .d(
        \sig_prgm_register/or_signal [620]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[620]) );
  d_ff \sig_prgm_register/genblk1[619].single_DFF  ( .d(
        \sig_prgm_register/or_signal [619]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[619]) );
  d_ff \sig_prgm_register/genblk1[618].single_DFF  ( .d(
        \sig_prgm_register/or_signal [618]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[618]) );
  d_ff \sig_prgm_register/genblk1[617].single_DFF  ( .d(
        \sig_prgm_register/or_signal [617]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[617]) );
  d_ff \sig_prgm_register/genblk1[616].single_DFF  ( .d(
        \sig_prgm_register/or_signal [616]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[616]) );
  d_ff \sig_prgm_register/genblk1[615].single_DFF  ( .d(
        \sig_prgm_register/or_signal [615]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[615]) );
  d_ff \sig_prgm_register/genblk1[614].single_DFF  ( .d(
        \sig_prgm_register/or_signal [614]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[614]) );
  d_ff \sig_prgm_register/genblk1[613].single_DFF  ( .d(
        \sig_prgm_register/or_signal [613]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[613]) );
  d_ff \sig_prgm_register/genblk1[612].single_DFF  ( .d(
        \sig_prgm_register/or_signal [612]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[612]) );
  d_ff \sig_prgm_register/genblk1[611].single_DFF  ( .d(
        \sig_prgm_register/or_signal [611]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[611]) );
  d_ff \sig_prgm_register/genblk1[610].single_DFF  ( .d(
        \sig_prgm_register/or_signal [610]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[610]) );
  d_ff \sig_prgm_register/genblk1[609].single_DFF  ( .d(
        \sig_prgm_register/or_signal [609]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[609]) );
  d_ff \sig_prgm_register/genblk1[608].single_DFF  ( .d(
        \sig_prgm_register/or_signal [608]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[608]) );
  d_ff \sig_prgm_register/genblk1[607].single_DFF  ( .d(
        \sig_prgm_register/or_signal [607]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[607]) );
  d_ff \sig_prgm_register/genblk1[606].single_DFF  ( .d(
        \sig_prgm_register/or_signal [606]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[606]) );
  d_ff \sig_prgm_register/genblk1[605].single_DFF  ( .d(
        \sig_prgm_register/or_signal [605]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[605]) );
  d_ff \sig_prgm_register/genblk1[604].single_DFF  ( .d(
        \sig_prgm_register/or_signal [604]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[604]) );
  d_ff \sig_prgm_register/genblk1[603].single_DFF  ( .d(
        \sig_prgm_register/or_signal [603]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[603]) );
  d_ff \sig_prgm_register/genblk1[602].single_DFF  ( .d(
        \sig_prgm_register/or_signal [602]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[602]) );
  d_ff \sig_prgm_register/genblk1[601].single_DFF  ( .d(
        \sig_prgm_register/or_signal [601]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[601]) );
  d_ff \sig_prgm_register/genblk1[600].single_DFF  ( .d(
        \sig_prgm_register/or_signal [600]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[600]) );
  d_ff \sig_prgm_register/genblk1[599].single_DFF  ( .d(
        \sig_prgm_register/or_signal [599]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[599]) );
  d_ff \sig_prgm_register/genblk1[598].single_DFF  ( .d(
        \sig_prgm_register/or_signal [598]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[598]) );
  d_ff \sig_prgm_register/genblk1[597].single_DFF  ( .d(
        \sig_prgm_register/or_signal [597]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[597]) );
  d_ff \sig_prgm_register/genblk1[596].single_DFF  ( .d(
        \sig_prgm_register/or_signal [596]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[596]) );
  d_ff \sig_prgm_register/genblk1[595].single_DFF  ( .d(
        \sig_prgm_register/or_signal [595]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[595]) );
  d_ff \sig_prgm_register/genblk1[594].single_DFF  ( .d(
        \sig_prgm_register/or_signal [594]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[594]) );
  d_ff \sig_prgm_register/genblk1[593].single_DFF  ( .d(
        \sig_prgm_register/or_signal [593]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[593]) );
  d_ff \sig_prgm_register/genblk1[592].single_DFF  ( .d(
        \sig_prgm_register/or_signal [592]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[592]) );
  d_ff \sig_prgm_register/genblk1[591].single_DFF  ( .d(
        \sig_prgm_register/or_signal [591]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[591]) );
  d_ff \sig_prgm_register/genblk1[590].single_DFF  ( .d(
        \sig_prgm_register/or_signal [590]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[590]) );
  d_ff \sig_prgm_register/genblk1[589].single_DFF  ( .d(
        \sig_prgm_register/or_signal [589]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[589]) );
  d_ff \sig_prgm_register/genblk1[588].single_DFF  ( .d(
        \sig_prgm_register/or_signal [588]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[588]) );
  d_ff \sig_prgm_register/genblk1[587].single_DFF  ( .d(
        \sig_prgm_register/or_signal [587]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[587]) );
  d_ff \sig_prgm_register/genblk1[586].single_DFF  ( .d(
        \sig_prgm_register/or_signal [586]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[586]) );
  d_ff \sig_prgm_register/genblk1[585].single_DFF  ( .d(
        \sig_prgm_register/or_signal [585]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[585]) );
  d_ff \sig_prgm_register/genblk1[584].single_DFF  ( .d(
        \sig_prgm_register/or_signal [584]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[584]) );
  d_ff \sig_prgm_register/genblk1[583].single_DFF  ( .d(
        \sig_prgm_register/or_signal [583]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[583]) );
  d_ff \sig_prgm_register/genblk1[582].single_DFF  ( .d(
        \sig_prgm_register/or_signal [582]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[582]) );
  d_ff \sig_prgm_register/genblk1[581].single_DFF  ( .d(
        \sig_prgm_register/or_signal [581]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[581]) );
  d_ff \sig_prgm_register/genblk1[580].single_DFF  ( .d(
        \sig_prgm_register/or_signal [580]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[580]) );
  d_ff \sig_prgm_register/genblk1[579].single_DFF  ( .d(
        \sig_prgm_register/or_signal [579]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[579]) );
  d_ff \sig_prgm_register/genblk1[578].single_DFF  ( .d(
        \sig_prgm_register/or_signal [578]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[578]) );
  d_ff \sig_prgm_register/genblk1[577].single_DFF  ( .d(
        \sig_prgm_register/or_signal [577]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[577]) );
  d_ff \sig_prgm_register/genblk1[576].single_DFF  ( .d(
        \sig_prgm_register/or_signal [576]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[576]) );
  d_ff \sig_prgm_register/genblk1[575].single_DFF  ( .d(
        \sig_prgm_register/or_signal [575]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[575]) );
  d_ff \sig_prgm_register/genblk1[574].single_DFF  ( .d(
        \sig_prgm_register/or_signal [574]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[574]) );
  d_ff \sig_prgm_register/genblk1[573].single_DFF  ( .d(
        \sig_prgm_register/or_signal [573]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[573]) );
  d_ff \sig_prgm_register/genblk1[572].single_DFF  ( .d(
        \sig_prgm_register/or_signal [572]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[572]) );
  d_ff \sig_prgm_register/genblk1[571].single_DFF  ( .d(
        \sig_prgm_register/or_signal [571]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[571]) );
  d_ff \sig_prgm_register/genblk1[570].single_DFF  ( .d(
        \sig_prgm_register/or_signal [570]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[570]) );
  d_ff \sig_prgm_register/genblk1[569].single_DFF  ( .d(
        \sig_prgm_register/or_signal [569]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[569]) );
  d_ff \sig_prgm_register/genblk1[568].single_DFF  ( .d(
        \sig_prgm_register/or_signal [568]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[568]) );
  d_ff \sig_prgm_register/genblk1[567].single_DFF  ( .d(
        \sig_prgm_register/or_signal [567]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[567]) );
  d_ff \sig_prgm_register/genblk1[566].single_DFF  ( .d(
        \sig_prgm_register/or_signal [566]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[566]) );
  d_ff \sig_prgm_register/genblk1[565].single_DFF  ( .d(
        \sig_prgm_register/or_signal [565]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[565]) );
  d_ff \sig_prgm_register/genblk1[564].single_DFF  ( .d(
        \sig_prgm_register/or_signal [564]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[564]) );
  d_ff \sig_prgm_register/genblk1[563].single_DFF  ( .d(
        \sig_prgm_register/or_signal [563]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[563]) );
  d_ff \sig_prgm_register/genblk1[562].single_DFF  ( .d(
        \sig_prgm_register/or_signal [562]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[562]) );
  d_ff \sig_prgm_register/genblk1[561].single_DFF  ( .d(
        \sig_prgm_register/or_signal [561]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[561]) );
  d_ff \sig_prgm_register/genblk1[560].single_DFF  ( .d(
        \sig_prgm_register/or_signal [560]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[560]) );
  d_ff \sig_prgm_register/genblk1[559].single_DFF  ( .d(
        \sig_prgm_register/or_signal [559]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[559]) );
  d_ff \sig_prgm_register/genblk1[558].single_DFF  ( .d(
        \sig_prgm_register/or_signal [558]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[558]) );
  d_ff \sig_prgm_register/genblk1[557].single_DFF  ( .d(
        \sig_prgm_register/or_signal [557]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[557]) );
  d_ff \sig_prgm_register/genblk1[556].single_DFF  ( .d(
        \sig_prgm_register/or_signal [556]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[556]) );
  d_ff \sig_prgm_register/genblk1[555].single_DFF  ( .d(
        \sig_prgm_register/or_signal [555]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[555]) );
  d_ff \sig_prgm_register/genblk1[554].single_DFF  ( .d(
        \sig_prgm_register/or_signal [554]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[554]) );
  d_ff \sig_prgm_register/genblk1[553].single_DFF  ( .d(
        \sig_prgm_register/or_signal [553]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[553]) );
  d_ff \sig_prgm_register/genblk1[552].single_DFF  ( .d(
        \sig_prgm_register/or_signal [552]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[552]) );
  d_ff \sig_prgm_register/genblk1[551].single_DFF  ( .d(
        \sig_prgm_register/or_signal [551]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[551]) );
  d_ff \sig_prgm_register/genblk1[550].single_DFF  ( .d(
        \sig_prgm_register/or_signal [550]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[550]) );
  d_ff \sig_prgm_register/genblk1[549].single_DFF  ( .d(
        \sig_prgm_register/or_signal [549]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[549]) );
  d_ff \sig_prgm_register/genblk1[548].single_DFF  ( .d(
        \sig_prgm_register/or_signal [548]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[548]) );
  d_ff \sig_prgm_register/genblk1[547].single_DFF  ( .d(
        \sig_prgm_register/or_signal [547]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[547]) );
  d_ff \sig_prgm_register/genblk1[546].single_DFF  ( .d(
        \sig_prgm_register/or_signal [546]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[546]) );
  d_ff \sig_prgm_register/genblk1[545].single_DFF  ( .d(
        \sig_prgm_register/or_signal [545]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[545]) );
  d_ff \sig_prgm_register/genblk1[544].single_DFF  ( .d(
        \sig_prgm_register/or_signal [544]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[544]) );
  d_ff \sig_prgm_register/genblk1[543].single_DFF  ( .d(
        \sig_prgm_register/or_signal [543]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[543]) );
  d_ff \sig_prgm_register/genblk1[542].single_DFF  ( .d(
        \sig_prgm_register/or_signal [542]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[542]) );
  d_ff \sig_prgm_register/genblk1[541].single_DFF  ( .d(
        \sig_prgm_register/or_signal [541]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[541]) );
  d_ff \sig_prgm_register/genblk1[540].single_DFF  ( .d(
        \sig_prgm_register/or_signal [540]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[540]) );
  d_ff \sig_prgm_register/genblk1[539].single_DFF  ( .d(
        \sig_prgm_register/or_signal [539]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[539]) );
  d_ff \sig_prgm_register/genblk1[538].single_DFF  ( .d(
        \sig_prgm_register/or_signal [538]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[538]) );
  d_ff \sig_prgm_register/genblk1[537].single_DFF  ( .d(
        \sig_prgm_register/or_signal [537]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[537]) );
  d_ff \sig_prgm_register/genblk1[536].single_DFF  ( .d(
        \sig_prgm_register/or_signal [536]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[536]) );
  d_ff \sig_prgm_register/genblk1[535].single_DFF  ( .d(
        \sig_prgm_register/or_signal [535]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[535]) );
  d_ff \sig_prgm_register/genblk1[534].single_DFF  ( .d(
        \sig_prgm_register/or_signal [534]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[534]) );
  d_ff \sig_prgm_register/genblk1[533].single_DFF  ( .d(
        \sig_prgm_register/or_signal [533]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[533]) );
  d_ff \sig_prgm_register/genblk1[532].single_DFF  ( .d(
        \sig_prgm_register/or_signal [532]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[532]) );
  d_ff \sig_prgm_register/genblk1[531].single_DFF  ( .d(
        \sig_prgm_register/or_signal [531]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[531]) );
  d_ff \sig_prgm_register/genblk1[530].single_DFF  ( .d(
        \sig_prgm_register/or_signal [530]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[530]) );
  d_ff \sig_prgm_register/genblk1[529].single_DFF  ( .d(
        \sig_prgm_register/or_signal [529]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[529]) );
  d_ff \sig_prgm_register/genblk1[528].single_DFF  ( .d(
        \sig_prgm_register/or_signal [528]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[528]) );
  d_ff \sig_prgm_register/genblk1[527].single_DFF  ( .d(
        \sig_prgm_register/or_signal [527]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[527]) );
  d_ff \sig_prgm_register/genblk1[526].single_DFF  ( .d(
        \sig_prgm_register/or_signal [526]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[526]) );
  d_ff \sig_prgm_register/genblk1[525].single_DFF  ( .d(
        \sig_prgm_register/or_signal [525]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[525]) );
  d_ff \sig_prgm_register/genblk1[524].single_DFF  ( .d(
        \sig_prgm_register/or_signal [524]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[524]) );
  d_ff \sig_prgm_register/genblk1[523].single_DFF  ( .d(
        \sig_prgm_register/or_signal [523]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[523]) );
  d_ff \sig_prgm_register/genblk1[522].single_DFF  ( .d(
        \sig_prgm_register/or_signal [522]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[522]) );
  d_ff \sig_prgm_register/genblk1[521].single_DFF  ( .d(
        \sig_prgm_register/or_signal [521]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[521]) );
  d_ff \sig_prgm_register/genblk1[520].single_DFF  ( .d(
        \sig_prgm_register/or_signal [520]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[520]) );
  d_ff \sig_prgm_register/genblk1[519].single_DFF  ( .d(
        \sig_prgm_register/or_signal [519]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[519]) );
  d_ff \sig_prgm_register/genblk1[518].single_DFF  ( .d(
        \sig_prgm_register/or_signal [518]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[518]) );
  d_ff \sig_prgm_register/genblk1[517].single_DFF  ( .d(
        \sig_prgm_register/or_signal [517]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[517]) );
  d_ff \sig_prgm_register/genblk1[516].single_DFF  ( .d(
        \sig_prgm_register/or_signal [516]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[516]) );
  d_ff \sig_prgm_register/genblk1[515].single_DFF  ( .d(
        \sig_prgm_register/or_signal [515]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[515]) );
  d_ff \sig_prgm_register/genblk1[514].single_DFF  ( .d(
        \sig_prgm_register/or_signal [514]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[514]) );
  d_ff \sig_prgm_register/genblk1[513].single_DFF  ( .d(
        \sig_prgm_register/or_signal [513]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[513]) );
  d_ff \sig_prgm_register/genblk1[512].single_DFF  ( .d(
        \sig_prgm_register/or_signal [512]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[512]) );
  d_ff \sig_prgm_register/genblk1[511].single_DFF  ( .d(
        \sig_prgm_register/or_signal [511]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[511]) );
  d_ff \sig_prgm_register/genblk1[510].single_DFF  ( .d(
        \sig_prgm_register/or_signal [510]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[510]) );
  d_ff \sig_prgm_register/genblk1[509].single_DFF  ( .d(
        \sig_prgm_register/or_signal [509]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[509]) );
  d_ff \sig_prgm_register/genblk1[508].single_DFF  ( .d(
        \sig_prgm_register/or_signal [508]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[508]) );
  d_ff \sig_prgm_register/genblk1[507].single_DFF  ( .d(
        \sig_prgm_register/or_signal [507]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[507]) );
  d_ff \sig_prgm_register/genblk1[506].single_DFF  ( .d(
        \sig_prgm_register/or_signal [506]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[506]) );
  d_ff \sig_prgm_register/genblk1[505].single_DFF  ( .d(
        \sig_prgm_register/or_signal [505]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[505]) );
  d_ff \sig_prgm_register/genblk1[504].single_DFF  ( .d(
        \sig_prgm_register/or_signal [504]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[504]) );
  d_ff \sig_prgm_register/genblk1[503].single_DFF  ( .d(
        \sig_prgm_register/or_signal [503]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[503]) );
  d_ff \sig_prgm_register/genblk1[502].single_DFF  ( .d(
        \sig_prgm_register/or_signal [502]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[502]) );
  d_ff \sig_prgm_register/genblk1[501].single_DFF  ( .d(
        \sig_prgm_register/or_signal [501]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[501]) );
  d_ff \sig_prgm_register/genblk1[500].single_DFF  ( .d(
        \sig_prgm_register/or_signal [500]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[500]) );
  d_ff \sig_prgm_register/genblk1[499].single_DFF  ( .d(
        \sig_prgm_register/or_signal [499]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[499]) );
  d_ff \sig_prgm_register/genblk1[498].single_DFF  ( .d(
        \sig_prgm_register/or_signal [498]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[498]) );
  d_ff \sig_prgm_register/genblk1[497].single_DFF  ( .d(
        \sig_prgm_register/or_signal [497]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[497]) );
  d_ff \sig_prgm_register/genblk1[496].single_DFF  ( .d(
        \sig_prgm_register/or_signal [496]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[496]) );
  d_ff \sig_prgm_register/genblk1[495].single_DFF  ( .d(
        \sig_prgm_register/or_signal [495]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[495]) );
  d_ff \sig_prgm_register/genblk1[494].single_DFF  ( .d(
        \sig_prgm_register/or_signal [494]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[494]) );
  d_ff \sig_prgm_register/genblk1[493].single_DFF  ( .d(
        \sig_prgm_register/or_signal [493]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[493]) );
  d_ff \sig_prgm_register/genblk1[492].single_DFF  ( .d(
        \sig_prgm_register/or_signal [492]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[492]) );
  d_ff \sig_prgm_register/genblk1[491].single_DFF  ( .d(
        \sig_prgm_register/or_signal [491]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[491]) );
  d_ff \sig_prgm_register/genblk1[490].single_DFF  ( .d(
        \sig_prgm_register/or_signal [490]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[490]) );
  d_ff \sig_prgm_register/genblk1[489].single_DFF  ( .d(
        \sig_prgm_register/or_signal [489]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[489]) );
  d_ff \sig_prgm_register/genblk1[488].single_DFF  ( .d(
        \sig_prgm_register/or_signal [488]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[488]) );
  d_ff \sig_prgm_register/genblk1[487].single_DFF  ( .d(
        \sig_prgm_register/or_signal [487]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[487]) );
  d_ff \sig_prgm_register/genblk1[486].single_DFF  ( .d(
        \sig_prgm_register/or_signal [486]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[486]) );
  d_ff \sig_prgm_register/genblk1[485].single_DFF  ( .d(
        \sig_prgm_register/or_signal [485]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[485]) );
  d_ff \sig_prgm_register/genblk1[484].single_DFF  ( .d(
        \sig_prgm_register/or_signal [484]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[484]) );
  d_ff \sig_prgm_register/genblk1[483].single_DFF  ( .d(
        \sig_prgm_register/or_signal [483]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[483]) );
  d_ff \sig_prgm_register/genblk1[482].single_DFF  ( .d(
        \sig_prgm_register/or_signal [482]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[482]) );
  d_ff \sig_prgm_register/genblk1[481].single_DFF  ( .d(
        \sig_prgm_register/or_signal [481]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[481]) );
  d_ff \sig_prgm_register/genblk1[480].single_DFF  ( .d(
        \sig_prgm_register/or_signal [480]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[480]) );
  d_ff \sig_prgm_register/genblk1[479].single_DFF  ( .d(
        \sig_prgm_register/or_signal [479]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[479]) );
  d_ff \sig_prgm_register/genblk1[478].single_DFF  ( .d(
        \sig_prgm_register/or_signal [478]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[478]) );
  d_ff \sig_prgm_register/genblk1[477].single_DFF  ( .d(
        \sig_prgm_register/or_signal [477]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[477]) );
  d_ff \sig_prgm_register/genblk1[476].single_DFF  ( .d(
        \sig_prgm_register/or_signal [476]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[476]) );
  d_ff \sig_prgm_register/genblk1[475].single_DFF  ( .d(
        \sig_prgm_register/or_signal [475]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[475]) );
  d_ff \sig_prgm_register/genblk1[474].single_DFF  ( .d(
        \sig_prgm_register/or_signal [474]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[474]) );
  d_ff \sig_prgm_register/genblk1[473].single_DFF  ( .d(
        \sig_prgm_register/or_signal [473]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[473]) );
  d_ff \sig_prgm_register/genblk1[472].single_DFF  ( .d(
        \sig_prgm_register/or_signal [472]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[472]) );
  d_ff \sig_prgm_register/genblk1[471].single_DFF  ( .d(
        \sig_prgm_register/or_signal [471]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[471]) );
  d_ff \sig_prgm_register/genblk1[470].single_DFF  ( .d(
        \sig_prgm_register/or_signal [470]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[470]) );
  d_ff \sig_prgm_register/genblk1[469].single_DFF  ( .d(
        \sig_prgm_register/or_signal [469]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[469]) );
  d_ff \sig_prgm_register/genblk1[468].single_DFF  ( .d(
        \sig_prgm_register/or_signal [468]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[468]) );
  d_ff \sig_prgm_register/genblk1[467].single_DFF  ( .d(
        \sig_prgm_register/or_signal [467]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[467]) );
  d_ff \sig_prgm_register/genblk1[466].single_DFF  ( .d(
        \sig_prgm_register/or_signal [466]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[466]) );
  d_ff \sig_prgm_register/genblk1[465].single_DFF  ( .d(
        \sig_prgm_register/or_signal [465]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[465]) );
  d_ff \sig_prgm_register/genblk1[464].single_DFF  ( .d(
        \sig_prgm_register/or_signal [464]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[464]) );
  d_ff \sig_prgm_register/genblk1[463].single_DFF  ( .d(
        \sig_prgm_register/or_signal [463]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[463]) );
  d_ff \sig_prgm_register/genblk1[462].single_DFF  ( .d(
        \sig_prgm_register/or_signal [462]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[462]) );
  d_ff \sig_prgm_register/genblk1[461].single_DFF  ( .d(
        \sig_prgm_register/or_signal [461]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[461]) );
  d_ff \sig_prgm_register/genblk1[460].single_DFF  ( .d(
        \sig_prgm_register/or_signal [460]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[460]) );
  d_ff \sig_prgm_register/genblk1[459].single_DFF  ( .d(
        \sig_prgm_register/or_signal [459]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[459]) );
  d_ff \sig_prgm_register/genblk1[458].single_DFF  ( .d(
        \sig_prgm_register/or_signal [458]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[458]) );
  d_ff \sig_prgm_register/genblk1[457].single_DFF  ( .d(
        \sig_prgm_register/or_signal [457]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[457]) );
  d_ff \sig_prgm_register/genblk1[456].single_DFF  ( .d(
        \sig_prgm_register/or_signal [456]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[456]) );
  d_ff \sig_prgm_register/genblk1[455].single_DFF  ( .d(
        \sig_prgm_register/or_signal [455]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[455]) );
  d_ff \sig_prgm_register/genblk1[454].single_DFF  ( .d(
        \sig_prgm_register/or_signal [454]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[454]) );
  d_ff \sig_prgm_register/genblk1[453].single_DFF  ( .d(
        \sig_prgm_register/or_signal [453]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[453]) );
  d_ff \sig_prgm_register/genblk1[452].single_DFF  ( .d(
        \sig_prgm_register/or_signal [452]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[452]) );
  d_ff \sig_prgm_register/genblk1[451].single_DFF  ( .d(
        \sig_prgm_register/or_signal [451]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[451]) );
  d_ff \sig_prgm_register/genblk1[450].single_DFF  ( .d(
        \sig_prgm_register/or_signal [450]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[450]) );
  d_ff \sig_prgm_register/genblk1[449].single_DFF  ( .d(
        \sig_prgm_register/or_signal [449]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[449]) );
  d_ff \sig_prgm_register/genblk1[448].single_DFF  ( .d(
        \sig_prgm_register/or_signal [448]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[448]) );
  d_ff \sig_prgm_register/genblk1[447].single_DFF  ( .d(
        \sig_prgm_register/or_signal [447]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[447]) );
  d_ff \sig_prgm_register/genblk1[446].single_DFF  ( .d(
        \sig_prgm_register/or_signal [446]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[446]) );
  d_ff \sig_prgm_register/genblk1[445].single_DFF  ( .d(
        \sig_prgm_register/or_signal [445]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[445]) );
  d_ff \sig_prgm_register/genblk1[444].single_DFF  ( .d(
        \sig_prgm_register/or_signal [444]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[444]) );
  d_ff \sig_prgm_register/genblk1[443].single_DFF  ( .d(
        \sig_prgm_register/or_signal [443]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[443]) );
  d_ff \sig_prgm_register/genblk1[442].single_DFF  ( .d(
        \sig_prgm_register/or_signal [442]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[442]) );
  d_ff \sig_prgm_register/genblk1[441].single_DFF  ( .d(
        \sig_prgm_register/or_signal [441]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[441]) );
  d_ff \sig_prgm_register/genblk1[440].single_DFF  ( .d(
        \sig_prgm_register/or_signal [440]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[440]) );
  d_ff \sig_prgm_register/genblk1[439].single_DFF  ( .d(
        \sig_prgm_register/or_signal [439]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[439]) );
  d_ff \sig_prgm_register/genblk1[438].single_DFF  ( .d(
        \sig_prgm_register/or_signal [438]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[438]) );
  d_ff \sig_prgm_register/genblk1[437].single_DFF  ( .d(
        \sig_prgm_register/or_signal [437]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[437]) );
  d_ff \sig_prgm_register/genblk1[436].single_DFF  ( .d(
        \sig_prgm_register/or_signal [436]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[436]) );
  d_ff \sig_prgm_register/genblk1[435].single_DFF  ( .d(
        \sig_prgm_register/or_signal [435]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[435]) );
  d_ff \sig_prgm_register/genblk1[434].single_DFF  ( .d(
        \sig_prgm_register/or_signal [434]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[434]) );
  d_ff \sig_prgm_register/genblk1[433].single_DFF  ( .d(
        \sig_prgm_register/or_signal [433]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[433]) );
  d_ff \sig_prgm_register/genblk1[432].single_DFF  ( .d(
        \sig_prgm_register/or_signal [432]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[432]) );
  d_ff \sig_prgm_register/genblk1[431].single_DFF  ( .d(
        \sig_prgm_register/or_signal [431]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[431]) );
  d_ff \sig_prgm_register/genblk1[430].single_DFF  ( .d(
        \sig_prgm_register/or_signal [430]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[430]) );
  d_ff \sig_prgm_register/genblk1[429].single_DFF  ( .d(
        \sig_prgm_register/or_signal [429]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[429]) );
  d_ff \sig_prgm_register/genblk1[428].single_DFF  ( .d(
        \sig_prgm_register/or_signal [428]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[428]) );
  d_ff \sig_prgm_register/genblk1[427].single_DFF  ( .d(
        \sig_prgm_register/or_signal [427]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[427]) );
  d_ff \sig_prgm_register/genblk1[426].single_DFF  ( .d(
        \sig_prgm_register/or_signal [426]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[426]) );
  d_ff \sig_prgm_register/genblk1[425].single_DFF  ( .d(
        \sig_prgm_register/or_signal [425]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[425]) );
  d_ff \sig_prgm_register/genblk1[424].single_DFF  ( .d(
        \sig_prgm_register/or_signal [424]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[424]) );
  d_ff \sig_prgm_register/genblk1[423].single_DFF  ( .d(
        \sig_prgm_register/or_signal [423]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[423]) );
  d_ff \sig_prgm_register/genblk1[422].single_DFF  ( .d(
        \sig_prgm_register/or_signal [422]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[422]) );
  d_ff \sig_prgm_register/genblk1[421].single_DFF  ( .d(
        \sig_prgm_register/or_signal [421]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[421]) );
  d_ff \sig_prgm_register/genblk1[420].single_DFF  ( .d(
        \sig_prgm_register/or_signal [420]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[420]) );
  d_ff \sig_prgm_register/genblk1[419].single_DFF  ( .d(
        \sig_prgm_register/or_signal [419]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[419]) );
  d_ff \sig_prgm_register/genblk1[418].single_DFF  ( .d(
        \sig_prgm_register/or_signal [418]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[418]) );
  d_ff \sig_prgm_register/genblk1[417].single_DFF  ( .d(
        \sig_prgm_register/or_signal [417]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[417]) );
  d_ff \sig_prgm_register/genblk1[416].single_DFF  ( .d(
        \sig_prgm_register/or_signal [416]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[416]) );
  d_ff \sig_prgm_register/genblk1[415].single_DFF  ( .d(
        \sig_prgm_register/or_signal [415]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[415]) );
  d_ff \sig_prgm_register/genblk1[414].single_DFF  ( .d(
        \sig_prgm_register/or_signal [414]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[414]) );
  d_ff \sig_prgm_register/genblk1[413].single_DFF  ( .d(
        \sig_prgm_register/or_signal [413]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[413]) );
  d_ff \sig_prgm_register/genblk1[412].single_DFF  ( .d(
        \sig_prgm_register/or_signal [412]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[412]) );
  d_ff \sig_prgm_register/genblk1[411].single_DFF  ( .d(
        \sig_prgm_register/or_signal [411]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[411]) );
  d_ff \sig_prgm_register/genblk1[410].single_DFF  ( .d(
        \sig_prgm_register/or_signal [410]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[410]) );
  d_ff \sig_prgm_register/genblk1[409].single_DFF  ( .d(
        \sig_prgm_register/or_signal [409]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[409]) );
  d_ff \sig_prgm_register/genblk1[408].single_DFF  ( .d(
        \sig_prgm_register/or_signal [408]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[408]) );
  d_ff \sig_prgm_register/genblk1[407].single_DFF  ( .d(
        \sig_prgm_register/or_signal [407]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[407]) );
  d_ff \sig_prgm_register/genblk1[406].single_DFF  ( .d(
        \sig_prgm_register/or_signal [406]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[406]) );
  d_ff \sig_prgm_register/genblk1[405].single_DFF  ( .d(
        \sig_prgm_register/or_signal [405]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[405]) );
  d_ff \sig_prgm_register/genblk1[404].single_DFF  ( .d(
        \sig_prgm_register/or_signal [404]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[404]) );
  d_ff \sig_prgm_register/genblk1[403].single_DFF  ( .d(
        \sig_prgm_register/or_signal [403]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[403]) );
  d_ff \sig_prgm_register/genblk1[402].single_DFF  ( .d(
        \sig_prgm_register/or_signal [402]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[402]) );
  d_ff \sig_prgm_register/genblk1[401].single_DFF  ( .d(
        \sig_prgm_register/or_signal [401]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[401]) );
  d_ff \sig_prgm_register/genblk1[400].single_DFF  ( .d(
        \sig_prgm_register/or_signal [400]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[400]) );
  d_ff \sig_prgm_register/genblk1[399].single_DFF  ( .d(
        \sig_prgm_register/or_signal [399]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[399]) );
  d_ff \sig_prgm_register/genblk1[398].single_DFF  ( .d(
        \sig_prgm_register/or_signal [398]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[398]) );
  d_ff \sig_prgm_register/genblk1[397].single_DFF  ( .d(
        \sig_prgm_register/or_signal [397]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[397]) );
  d_ff \sig_prgm_register/genblk1[396].single_DFF  ( .d(
        \sig_prgm_register/or_signal [396]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[396]) );
  d_ff \sig_prgm_register/genblk1[395].single_DFF  ( .d(
        \sig_prgm_register/or_signal [395]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[395]) );
  d_ff \sig_prgm_register/genblk1[394].single_DFF  ( .d(
        \sig_prgm_register/or_signal [394]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[394]) );
  d_ff \sig_prgm_register/genblk1[393].single_DFF  ( .d(
        \sig_prgm_register/or_signal [393]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[393]) );
  d_ff \sig_prgm_register/genblk1[392].single_DFF  ( .d(
        \sig_prgm_register/or_signal [392]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[392]) );
  d_ff \sig_prgm_register/genblk1[391].single_DFF  ( .d(
        \sig_prgm_register/or_signal [391]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[391]) );
  d_ff \sig_prgm_register/genblk1[390].single_DFF  ( .d(
        \sig_prgm_register/or_signal [390]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[390]) );
  d_ff \sig_prgm_register/genblk1[389].single_DFF  ( .d(
        \sig_prgm_register/or_signal [389]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[389]) );
  d_ff \sig_prgm_register/genblk1[388].single_DFF  ( .d(
        \sig_prgm_register/or_signal [388]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[388]) );
  d_ff \sig_prgm_register/genblk1[387].single_DFF  ( .d(
        \sig_prgm_register/or_signal [387]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[387]) );
  d_ff \sig_prgm_register/genblk1[386].single_DFF  ( .d(
        \sig_prgm_register/or_signal [386]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[386]) );
  d_ff \sig_prgm_register/genblk1[385].single_DFF  ( .d(
        \sig_prgm_register/or_signal [385]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[385]) );
  d_ff \sig_prgm_register/genblk1[384].single_DFF  ( .d(
        \sig_prgm_register/or_signal [384]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[384]) );
  d_ff \sig_prgm_register/genblk1[383].single_DFF  ( .d(
        \sig_prgm_register/or_signal [383]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[383]) );
  d_ff \sig_prgm_register/genblk1[382].single_DFF  ( .d(
        \sig_prgm_register/or_signal [382]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[382]) );
  d_ff \sig_prgm_register/genblk1[381].single_DFF  ( .d(
        \sig_prgm_register/or_signal [381]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[381]) );
  d_ff \sig_prgm_register/genblk1[380].single_DFF  ( .d(
        \sig_prgm_register/or_signal [380]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[380]) );
  d_ff \sig_prgm_register/genblk1[379].single_DFF  ( .d(
        \sig_prgm_register/or_signal [379]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[379]) );
  d_ff \sig_prgm_register/genblk1[378].single_DFF  ( .d(
        \sig_prgm_register/or_signal [378]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[378]) );
  d_ff \sig_prgm_register/genblk1[377].single_DFF  ( .d(
        \sig_prgm_register/or_signal [377]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[377]) );
  d_ff \sig_prgm_register/genblk1[376].single_DFF  ( .d(
        \sig_prgm_register/or_signal [376]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[376]) );
  d_ff \sig_prgm_register/genblk1[375].single_DFF  ( .d(
        \sig_prgm_register/or_signal [375]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[375]) );
  d_ff \sig_prgm_register/genblk1[374].single_DFF  ( .d(
        \sig_prgm_register/or_signal [374]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[374]) );
  d_ff \sig_prgm_register/genblk1[373].single_DFF  ( .d(
        \sig_prgm_register/or_signal [373]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[373]) );
  d_ff \sig_prgm_register/genblk1[372].single_DFF  ( .d(
        \sig_prgm_register/or_signal [372]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[372]) );
  d_ff \sig_prgm_register/genblk1[371].single_DFF  ( .d(
        \sig_prgm_register/or_signal [371]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[371]) );
  d_ff \sig_prgm_register/genblk1[370].single_DFF  ( .d(
        \sig_prgm_register/or_signal [370]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[370]) );
  d_ff \sig_prgm_register/genblk1[369].single_DFF  ( .d(
        \sig_prgm_register/or_signal [369]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[369]) );
  d_ff \sig_prgm_register/genblk1[368].single_DFF  ( .d(
        \sig_prgm_register/or_signal [368]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[368]) );
  d_ff \sig_prgm_register/genblk1[367].single_DFF  ( .d(
        \sig_prgm_register/or_signal [367]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[367]) );
  d_ff \sig_prgm_register/genblk1[366].single_DFF  ( .d(
        \sig_prgm_register/or_signal [366]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[366]) );
  d_ff \sig_prgm_register/genblk1[365].single_DFF  ( .d(
        \sig_prgm_register/or_signal [365]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[365]) );
  d_ff \sig_prgm_register/genblk1[364].single_DFF  ( .d(
        \sig_prgm_register/or_signal [364]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[364]) );
  d_ff \sig_prgm_register/genblk1[363].single_DFF  ( .d(
        \sig_prgm_register/or_signal [363]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[363]) );
  d_ff \sig_prgm_register/genblk1[362].single_DFF  ( .d(
        \sig_prgm_register/or_signal [362]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[362]) );
  d_ff \sig_prgm_register/genblk1[361].single_DFF  ( .d(
        \sig_prgm_register/or_signal [361]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[361]) );
  d_ff \sig_prgm_register/genblk1[360].single_DFF  ( .d(
        \sig_prgm_register/or_signal [360]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[360]) );
  d_ff \sig_prgm_register/genblk1[359].single_DFF  ( .d(
        \sig_prgm_register/or_signal [359]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[359]) );
  d_ff \sig_prgm_register/genblk1[358].single_DFF  ( .d(
        \sig_prgm_register/or_signal [358]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[358]) );
  d_ff \sig_prgm_register/genblk1[357].single_DFF  ( .d(
        \sig_prgm_register/or_signal [357]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[357]) );
  d_ff \sig_prgm_register/genblk1[356].single_DFF  ( .d(
        \sig_prgm_register/or_signal [356]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[356]) );
  d_ff \sig_prgm_register/genblk1[355].single_DFF  ( .d(
        \sig_prgm_register/or_signal [355]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[355]) );
  d_ff \sig_prgm_register/genblk1[354].single_DFF  ( .d(
        \sig_prgm_register/or_signal [354]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[354]) );
  d_ff \sig_prgm_register/genblk1[353].single_DFF  ( .d(
        \sig_prgm_register/or_signal [353]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[353]) );
  d_ff \sig_prgm_register/genblk1[352].single_DFF  ( .d(
        \sig_prgm_register/or_signal [352]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[352]) );
  d_ff \sig_prgm_register/genblk1[351].single_DFF  ( .d(
        \sig_prgm_register/or_signal [351]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[351]) );
  d_ff \sig_prgm_register/genblk1[350].single_DFF  ( .d(
        \sig_prgm_register/or_signal [350]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[350]) );
  d_ff \sig_prgm_register/genblk1[349].single_DFF  ( .d(
        \sig_prgm_register/or_signal [349]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[349]) );
  d_ff \sig_prgm_register/genblk1[348].single_DFF  ( .d(
        \sig_prgm_register/or_signal [348]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[348]) );
  d_ff \sig_prgm_register/genblk1[347].single_DFF  ( .d(
        \sig_prgm_register/or_signal [347]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[347]) );
  d_ff \sig_prgm_register/genblk1[346].single_DFF  ( .d(
        \sig_prgm_register/or_signal [346]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[346]) );
  d_ff \sig_prgm_register/genblk1[345].single_DFF  ( .d(
        \sig_prgm_register/or_signal [345]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[345]) );
  d_ff \sig_prgm_register/genblk1[344].single_DFF  ( .d(
        \sig_prgm_register/or_signal [344]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[344]) );
  d_ff \sig_prgm_register/genblk1[343].single_DFF  ( .d(
        \sig_prgm_register/or_signal [343]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[343]) );
  d_ff \sig_prgm_register/genblk1[342].single_DFF  ( .d(
        \sig_prgm_register/or_signal [342]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[342]) );
  d_ff \sig_prgm_register/genblk1[341].single_DFF  ( .d(
        \sig_prgm_register/or_signal [341]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[341]) );
  d_ff \sig_prgm_register/genblk1[340].single_DFF  ( .d(
        \sig_prgm_register/or_signal [340]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[340]) );
  d_ff \sig_prgm_register/genblk1[339].single_DFF  ( .d(
        \sig_prgm_register/or_signal [339]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[339]) );
  d_ff \sig_prgm_register/genblk1[338].single_DFF  ( .d(
        \sig_prgm_register/or_signal [338]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[338]) );
  d_ff \sig_prgm_register/genblk1[337].single_DFF  ( .d(
        \sig_prgm_register/or_signal [337]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[337]) );
  d_ff \sig_prgm_register/genblk1[336].single_DFF  ( .d(
        \sig_prgm_register/or_signal [336]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[336]) );
  d_ff \sig_prgm_register/genblk1[335].single_DFF  ( .d(
        \sig_prgm_register/or_signal [335]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[335]) );
  d_ff \sig_prgm_register/genblk1[334].single_DFF  ( .d(
        \sig_prgm_register/or_signal [334]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[334]) );
  d_ff \sig_prgm_register/genblk1[333].single_DFF  ( .d(
        \sig_prgm_register/or_signal [333]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[333]) );
  d_ff \sig_prgm_register/genblk1[332].single_DFF  ( .d(
        \sig_prgm_register/or_signal [332]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[332]) );
  d_ff \sig_prgm_register/genblk1[331].single_DFF  ( .d(
        \sig_prgm_register/or_signal [331]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[331]) );
  d_ff \sig_prgm_register/genblk1[330].single_DFF  ( .d(
        \sig_prgm_register/or_signal [330]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[330]) );
  d_ff \sig_prgm_register/genblk1[329].single_DFF  ( .d(
        \sig_prgm_register/or_signal [329]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[329]) );
  d_ff \sig_prgm_register/genblk1[328].single_DFF  ( .d(
        \sig_prgm_register/or_signal [328]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[328]) );
  d_ff \sig_prgm_register/genblk1[327].single_DFF  ( .d(
        \sig_prgm_register/or_signal [327]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[327]) );
  d_ff \sig_prgm_register/genblk1[326].single_DFF  ( .d(
        \sig_prgm_register/or_signal [326]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[326]) );
  d_ff \sig_prgm_register/genblk1[325].single_DFF  ( .d(
        \sig_prgm_register/or_signal [325]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[325]) );
  d_ff \sig_prgm_register/genblk1[324].single_DFF  ( .d(
        \sig_prgm_register/or_signal [324]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[324]) );
  d_ff \sig_prgm_register/genblk1[323].single_DFF  ( .d(
        \sig_prgm_register/or_signal [323]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[323]) );
  d_ff \sig_prgm_register/genblk1[322].single_DFF  ( .d(
        \sig_prgm_register/or_signal [322]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[322]) );
  d_ff \sig_prgm_register/genblk1[321].single_DFF  ( .d(
        \sig_prgm_register/or_signal [321]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[321]) );
  d_ff \sig_prgm_register/genblk1[320].single_DFF  ( .d(
        \sig_prgm_register/or_signal [320]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[320]) );
  d_ff \sig_prgm_register/genblk1[319].single_DFF  ( .d(
        \sig_prgm_register/or_signal [319]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[319]) );
  d_ff \sig_prgm_register/genblk1[318].single_DFF  ( .d(
        \sig_prgm_register/or_signal [318]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[318]) );
  d_ff \sig_prgm_register/genblk1[317].single_DFF  ( .d(
        \sig_prgm_register/or_signal [317]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[317]) );
  d_ff \sig_prgm_register/genblk1[316].single_DFF  ( .d(
        \sig_prgm_register/or_signal [316]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[316]) );
  d_ff \sig_prgm_register/genblk1[315].single_DFF  ( .d(
        \sig_prgm_register/or_signal [315]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[315]) );
  d_ff \sig_prgm_register/genblk1[314].single_DFF  ( .d(
        \sig_prgm_register/or_signal [314]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[314]) );
  d_ff \sig_prgm_register/genblk1[313].single_DFF  ( .d(
        \sig_prgm_register/or_signal [313]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[313]) );
  d_ff \sig_prgm_register/genblk1[312].single_DFF  ( .d(
        \sig_prgm_register/or_signal [312]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[312]) );
  d_ff \sig_prgm_register/genblk1[311].single_DFF  ( .d(
        \sig_prgm_register/or_signal [311]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[311]) );
  d_ff \sig_prgm_register/genblk1[310].single_DFF  ( .d(
        \sig_prgm_register/or_signal [310]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[310]) );
  d_ff \sig_prgm_register/genblk1[309].single_DFF  ( .d(
        \sig_prgm_register/or_signal [309]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[309]) );
  d_ff \sig_prgm_register/genblk1[308].single_DFF  ( .d(
        \sig_prgm_register/or_signal [308]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[308]) );
  d_ff \sig_prgm_register/genblk1[307].single_DFF  ( .d(
        \sig_prgm_register/or_signal [307]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[307]) );
  d_ff \sig_prgm_register/genblk1[306].single_DFF  ( .d(
        \sig_prgm_register/or_signal [306]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[306]) );
  d_ff \sig_prgm_register/genblk1[305].single_DFF  ( .d(
        \sig_prgm_register/or_signal [305]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[305]) );
  d_ff \sig_prgm_register/genblk1[304].single_DFF  ( .d(
        \sig_prgm_register/or_signal [304]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[304]) );
  d_ff \sig_prgm_register/genblk1[303].single_DFF  ( .d(
        \sig_prgm_register/or_signal [303]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[303]) );
  d_ff \sig_prgm_register/genblk1[302].single_DFF  ( .d(
        \sig_prgm_register/or_signal [302]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[302]) );
  d_ff \sig_prgm_register/genblk1[301].single_DFF  ( .d(
        \sig_prgm_register/or_signal [301]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[301]) );
  d_ff \sig_prgm_register/genblk1[300].single_DFF  ( .d(
        \sig_prgm_register/or_signal [300]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[300]) );
  d_ff \sig_prgm_register/genblk1[299].single_DFF  ( .d(
        \sig_prgm_register/or_signal [299]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[299]) );
  d_ff \sig_prgm_register/genblk1[298].single_DFF  ( .d(
        \sig_prgm_register/or_signal [298]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[298]) );
  d_ff \sig_prgm_register/genblk1[297].single_DFF  ( .d(
        \sig_prgm_register/or_signal [297]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[297]) );
  d_ff \sig_prgm_register/genblk1[296].single_DFF  ( .d(
        \sig_prgm_register/or_signal [296]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[296]) );
  d_ff \sig_prgm_register/genblk1[295].single_DFF  ( .d(
        \sig_prgm_register/or_signal [295]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[295]) );
  d_ff \sig_prgm_register/genblk1[294].single_DFF  ( .d(
        \sig_prgm_register/or_signal [294]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[294]) );
  d_ff \sig_prgm_register/genblk1[293].single_DFF  ( .d(
        \sig_prgm_register/or_signal [293]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[293]) );
  d_ff \sig_prgm_register/genblk1[292].single_DFF  ( .d(
        \sig_prgm_register/or_signal [292]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[292]) );
  d_ff \sig_prgm_register/genblk1[291].single_DFF  ( .d(
        \sig_prgm_register/or_signal [291]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[291]) );
  d_ff \sig_prgm_register/genblk1[290].single_DFF  ( .d(
        \sig_prgm_register/or_signal [290]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[290]) );
  d_ff \sig_prgm_register/genblk1[289].single_DFF  ( .d(
        \sig_prgm_register/or_signal [289]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[289]) );
  d_ff \sig_prgm_register/genblk1[288].single_DFF  ( .d(
        \sig_prgm_register/or_signal [288]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[288]) );
  d_ff \sig_prgm_register/genblk1[287].single_DFF  ( .d(
        \sig_prgm_register/or_signal [287]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[287]) );
  d_ff \sig_prgm_register/genblk1[286].single_DFF  ( .d(
        \sig_prgm_register/or_signal [286]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[286]) );
  d_ff \sig_prgm_register/genblk1[285].single_DFF  ( .d(
        \sig_prgm_register/or_signal [285]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[285]) );
  d_ff \sig_prgm_register/genblk1[284].single_DFF  ( .d(
        \sig_prgm_register/or_signal [284]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[284]) );
  d_ff \sig_prgm_register/genblk1[283].single_DFF  ( .d(
        \sig_prgm_register/or_signal [283]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[283]) );
  d_ff \sig_prgm_register/genblk1[282].single_DFF  ( .d(
        \sig_prgm_register/or_signal [282]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[282]) );
  d_ff \sig_prgm_register/genblk1[281].single_DFF  ( .d(
        \sig_prgm_register/or_signal [281]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[281]) );
  d_ff \sig_prgm_register/genblk1[280].single_DFF  ( .d(
        \sig_prgm_register/or_signal [280]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[280]) );
  d_ff \sig_prgm_register/genblk1[279].single_DFF  ( .d(
        \sig_prgm_register/or_signal [279]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[279]) );
  d_ff \sig_prgm_register/genblk1[278].single_DFF  ( .d(
        \sig_prgm_register/or_signal [278]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[278]) );
  d_ff \sig_prgm_register/genblk1[277].single_DFF  ( .d(
        \sig_prgm_register/or_signal [277]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[277]) );
  d_ff \sig_prgm_register/genblk1[276].single_DFF  ( .d(
        \sig_prgm_register/or_signal [276]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[276]) );
  d_ff \sig_prgm_register/genblk1[275].single_DFF  ( .d(
        \sig_prgm_register/or_signal [275]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[275]) );
  d_ff \sig_prgm_register/genblk1[274].single_DFF  ( .d(
        \sig_prgm_register/or_signal [274]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[274]) );
  d_ff \sig_prgm_register/genblk1[273].single_DFF  ( .d(
        \sig_prgm_register/or_signal [273]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[273]) );
  d_ff \sig_prgm_register/genblk1[272].single_DFF  ( .d(
        \sig_prgm_register/or_signal [272]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[272]) );
  d_ff \sig_prgm_register/genblk1[271].single_DFF  ( .d(
        \sig_prgm_register/or_signal [271]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[271]) );
  d_ff \sig_prgm_register/genblk1[270].single_DFF  ( .d(
        \sig_prgm_register/or_signal [270]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[270]) );
  d_ff \sig_prgm_register/genblk1[269].single_DFF  ( .d(
        \sig_prgm_register/or_signal [269]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[269]) );
  d_ff \sig_prgm_register/genblk1[268].single_DFF  ( .d(
        \sig_prgm_register/or_signal [268]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[268]) );
  d_ff \sig_prgm_register/genblk1[267].single_DFF  ( .d(
        \sig_prgm_register/or_signal [267]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[267]) );
  d_ff \sig_prgm_register/genblk1[266].single_DFF  ( .d(
        \sig_prgm_register/or_signal [266]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[266]) );
  d_ff \sig_prgm_register/genblk1[265].single_DFF  ( .d(
        \sig_prgm_register/or_signal [265]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[265]) );
  d_ff \sig_prgm_register/genblk1[264].single_DFF  ( .d(
        \sig_prgm_register/or_signal [264]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[264]) );
  d_ff \sig_prgm_register/genblk1[263].single_DFF  ( .d(
        \sig_prgm_register/or_signal [263]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[263]) );
  d_ff \sig_prgm_register/genblk1[262].single_DFF  ( .d(
        \sig_prgm_register/or_signal [262]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[262]) );
  d_ff \sig_prgm_register/genblk1[261].single_DFF  ( .d(
        \sig_prgm_register/or_signal [261]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[261]) );
  d_ff \sig_prgm_register/genblk1[260].single_DFF  ( .d(
        \sig_prgm_register/or_signal [260]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[260]) );
  d_ff \sig_prgm_register/genblk1[259].single_DFF  ( .d(
        \sig_prgm_register/or_signal [259]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[259]) );
  d_ff \sig_prgm_register/genblk1[258].single_DFF  ( .d(
        \sig_prgm_register/or_signal [258]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[258]) );
  d_ff \sig_prgm_register/genblk1[257].single_DFF  ( .d(
        \sig_prgm_register/or_signal [257]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[257]) );
  d_ff \sig_prgm_register/genblk1[256].single_DFF  ( .d(
        \sig_prgm_register/or_signal [256]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[256]) );
  d_ff \sig_prgm_register/genblk1[255].single_DFF  ( .d(
        \sig_prgm_register/or_signal [255]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[255]) );
  d_ff \sig_prgm_register/genblk1[254].single_DFF  ( .d(
        \sig_prgm_register/or_signal [254]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[254]) );
  d_ff \sig_prgm_register/genblk1[253].single_DFF  ( .d(
        \sig_prgm_register/or_signal [253]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[253]) );
  d_ff \sig_prgm_register/genblk1[252].single_DFF  ( .d(
        \sig_prgm_register/or_signal [252]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[252]) );
  d_ff \sig_prgm_register/genblk1[251].single_DFF  ( .d(
        \sig_prgm_register/or_signal [251]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[251]) );
  d_ff \sig_prgm_register/genblk1[250].single_DFF  ( .d(
        \sig_prgm_register/or_signal [250]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[250]) );
  d_ff \sig_prgm_register/genblk1[249].single_DFF  ( .d(
        \sig_prgm_register/or_signal [249]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[249]) );
  d_ff \sig_prgm_register/genblk1[248].single_DFF  ( .d(
        \sig_prgm_register/or_signal [248]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[248]) );
  d_ff \sig_prgm_register/genblk1[247].single_DFF  ( .d(
        \sig_prgm_register/or_signal [247]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[247]) );
  d_ff \sig_prgm_register/genblk1[246].single_DFF  ( .d(
        \sig_prgm_register/or_signal [246]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[246]) );
  d_ff \sig_prgm_register/genblk1[245].single_DFF  ( .d(
        \sig_prgm_register/or_signal [245]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[245]) );
  d_ff \sig_prgm_register/genblk1[244].single_DFF  ( .d(
        \sig_prgm_register/or_signal [244]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[244]) );
  d_ff \sig_prgm_register/genblk1[243].single_DFF  ( .d(
        \sig_prgm_register/or_signal [243]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[243]) );
  d_ff \sig_prgm_register/genblk1[242].single_DFF  ( .d(
        \sig_prgm_register/or_signal [242]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[242]) );
  d_ff \sig_prgm_register/genblk1[241].single_DFF  ( .d(
        \sig_prgm_register/or_signal [241]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[241]) );
  d_ff \sig_prgm_register/genblk1[240].single_DFF  ( .d(
        \sig_prgm_register/or_signal [240]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[240]) );
  d_ff \sig_prgm_register/genblk1[239].single_DFF  ( .d(
        \sig_prgm_register/or_signal [239]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[239]) );
  d_ff \sig_prgm_register/genblk1[238].single_DFF  ( .d(
        \sig_prgm_register/or_signal [238]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[238]) );
  d_ff \sig_prgm_register/genblk1[237].single_DFF  ( .d(
        \sig_prgm_register/or_signal [237]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[237]) );
  d_ff \sig_prgm_register/genblk1[236].single_DFF  ( .d(
        \sig_prgm_register/or_signal [236]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[236]) );
  d_ff \sig_prgm_register/genblk1[235].single_DFF  ( .d(
        \sig_prgm_register/or_signal [235]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[235]) );
  d_ff \sig_prgm_register/genblk1[234].single_DFF  ( .d(
        \sig_prgm_register/or_signal [234]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[234]) );
  d_ff \sig_prgm_register/genblk1[233].single_DFF  ( .d(
        \sig_prgm_register/or_signal [233]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[233]) );
  d_ff \sig_prgm_register/genblk1[232].single_DFF  ( .d(
        \sig_prgm_register/or_signal [232]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[232]) );
  d_ff \sig_prgm_register/genblk1[231].single_DFF  ( .d(
        \sig_prgm_register/or_signal [231]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[231]) );
  d_ff \sig_prgm_register/genblk1[230].single_DFF  ( .d(
        \sig_prgm_register/or_signal [230]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[230]) );
  d_ff \sig_prgm_register/genblk1[229].single_DFF  ( .d(
        \sig_prgm_register/or_signal [229]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[229]) );
  d_ff \sig_prgm_register/genblk1[228].single_DFF  ( .d(
        \sig_prgm_register/or_signal [228]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[228]) );
  d_ff \sig_prgm_register/genblk1[227].single_DFF  ( .d(
        \sig_prgm_register/or_signal [227]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[227]) );
  d_ff \sig_prgm_register/genblk1[226].single_DFF  ( .d(
        \sig_prgm_register/or_signal [226]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[226]) );
  d_ff \sig_prgm_register/genblk1[225].single_DFF  ( .d(
        \sig_prgm_register/or_signal [225]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[225]) );
  d_ff \sig_prgm_register/genblk1[224].single_DFF  ( .d(
        \sig_prgm_register/or_signal [224]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[224]) );
  d_ff \sig_prgm_register/genblk1[223].single_DFF  ( .d(
        \sig_prgm_register/or_signal [223]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[223]) );
  d_ff \sig_prgm_register/genblk1[222].single_DFF  ( .d(
        \sig_prgm_register/or_signal [222]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[222]) );
  d_ff \sig_prgm_register/genblk1[221].single_DFF  ( .d(
        \sig_prgm_register/or_signal [221]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[221]) );
  d_ff \sig_prgm_register/genblk1[220].single_DFF  ( .d(
        \sig_prgm_register/or_signal [220]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[220]) );
  d_ff \sig_prgm_register/genblk1[219].single_DFF  ( .d(
        \sig_prgm_register/or_signal [219]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[219]) );
  d_ff \sig_prgm_register/genblk1[218].single_DFF  ( .d(
        \sig_prgm_register/or_signal [218]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[218]) );
  d_ff \sig_prgm_register/genblk1[217].single_DFF  ( .d(
        \sig_prgm_register/or_signal [217]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[217]) );
  d_ff \sig_prgm_register/genblk1[216].single_DFF  ( .d(
        \sig_prgm_register/or_signal [216]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[216]) );
  d_ff \sig_prgm_register/genblk1[215].single_DFF  ( .d(
        \sig_prgm_register/or_signal [215]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[215]) );
  d_ff \sig_prgm_register/genblk1[214].single_DFF  ( .d(
        \sig_prgm_register/or_signal [214]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[214]) );
  d_ff \sig_prgm_register/genblk1[213].single_DFF  ( .d(
        \sig_prgm_register/or_signal [213]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[213]) );
  d_ff \sig_prgm_register/genblk1[212].single_DFF  ( .d(
        \sig_prgm_register/or_signal [212]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[212]) );
  d_ff \sig_prgm_register/genblk1[211].single_DFF  ( .d(
        \sig_prgm_register/or_signal [211]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[211]) );
  d_ff \sig_prgm_register/genblk1[210].single_DFF  ( .d(
        \sig_prgm_register/or_signal [210]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[210]) );
  d_ff \sig_prgm_register/genblk1[209].single_DFF  ( .d(
        \sig_prgm_register/or_signal [209]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[209]) );
  d_ff \sig_prgm_register/genblk1[208].single_DFF  ( .d(
        \sig_prgm_register/or_signal [208]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[208]) );
  d_ff \sig_prgm_register/genblk1[207].single_DFF  ( .d(
        \sig_prgm_register/or_signal [207]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[207]) );
  d_ff \sig_prgm_register/genblk1[206].single_DFF  ( .d(
        \sig_prgm_register/or_signal [206]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[206]) );
  d_ff \sig_prgm_register/genblk1[205].single_DFF  ( .d(
        \sig_prgm_register/or_signal [205]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[205]) );
  d_ff \sig_prgm_register/genblk1[204].single_DFF  ( .d(
        \sig_prgm_register/or_signal [204]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[204]) );
  d_ff \sig_prgm_register/genblk1[203].single_DFF  ( .d(
        \sig_prgm_register/or_signal [203]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[203]) );
  d_ff \sig_prgm_register/genblk1[202].single_DFF  ( .d(
        \sig_prgm_register/or_signal [202]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[202]) );
  d_ff \sig_prgm_register/genblk1[201].single_DFF  ( .d(
        \sig_prgm_register/or_signal [201]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[201]) );
  d_ff \sig_prgm_register/genblk1[200].single_DFF  ( .d(
        \sig_prgm_register/or_signal [200]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[200]) );
  d_ff \sig_prgm_register/genblk1[199].single_DFF  ( .d(
        \sig_prgm_register/or_signal [199]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[199]) );
  d_ff \sig_prgm_register/genblk1[198].single_DFF  ( .d(
        \sig_prgm_register/or_signal [198]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[198]) );
  d_ff \sig_prgm_register/genblk1[197].single_DFF  ( .d(
        \sig_prgm_register/or_signal [197]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[197]) );
  d_ff \sig_prgm_register/genblk1[196].single_DFF  ( .d(
        \sig_prgm_register/or_signal [196]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[196]) );
  d_ff \sig_prgm_register/genblk1[195].single_DFF  ( .d(
        \sig_prgm_register/or_signal [195]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[195]) );
  d_ff \sig_prgm_register/genblk1[194].single_DFF  ( .d(
        \sig_prgm_register/or_signal [194]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[194]) );
  d_ff \sig_prgm_register/genblk1[193].single_DFF  ( .d(
        \sig_prgm_register/or_signal [193]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[193]) );
  d_ff \sig_prgm_register/genblk1[192].single_DFF  ( .d(
        \sig_prgm_register/or_signal [192]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[192]) );
  d_ff \sig_prgm_register/genblk1[191].single_DFF  ( .d(
        \sig_prgm_register/or_signal [191]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[191]) );
  d_ff \sig_prgm_register/genblk1[190].single_DFF  ( .d(
        \sig_prgm_register/or_signal [190]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[190]) );
  d_ff \sig_prgm_register/genblk1[189].single_DFF  ( .d(
        \sig_prgm_register/or_signal [189]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[189]) );
  d_ff \sig_prgm_register/genblk1[188].single_DFF  ( .d(
        \sig_prgm_register/or_signal [188]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[188]) );
  d_ff \sig_prgm_register/genblk1[187].single_DFF  ( .d(
        \sig_prgm_register/or_signal [187]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[187]) );
  d_ff \sig_prgm_register/genblk1[186].single_DFF  ( .d(
        \sig_prgm_register/or_signal [186]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[186]) );
  d_ff \sig_prgm_register/genblk1[185].single_DFF  ( .d(
        \sig_prgm_register/or_signal [185]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[185]) );
  d_ff \sig_prgm_register/genblk1[184].single_DFF  ( .d(
        \sig_prgm_register/or_signal [184]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[184]) );
  d_ff \sig_prgm_register/genblk1[183].single_DFF  ( .d(
        \sig_prgm_register/or_signal [183]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[183]) );
  d_ff \sig_prgm_register/genblk1[182].single_DFF  ( .d(
        \sig_prgm_register/or_signal [182]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[182]) );
  d_ff \sig_prgm_register/genblk1[181].single_DFF  ( .d(
        \sig_prgm_register/or_signal [181]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[181]) );
  d_ff \sig_prgm_register/genblk1[180].single_DFF  ( .d(
        \sig_prgm_register/or_signal [180]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[180]) );
  d_ff \sig_prgm_register/genblk1[179].single_DFF  ( .d(
        \sig_prgm_register/or_signal [179]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[179]) );
  d_ff \sig_prgm_register/genblk1[178].single_DFF  ( .d(
        \sig_prgm_register/or_signal [178]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[178]) );
  d_ff \sig_prgm_register/genblk1[177].single_DFF  ( .d(
        \sig_prgm_register/or_signal [177]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[177]) );
  d_ff \sig_prgm_register/genblk1[176].single_DFF  ( .d(
        \sig_prgm_register/or_signal [176]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[176]) );
  d_ff \sig_prgm_register/genblk1[175].single_DFF  ( .d(
        \sig_prgm_register/or_signal [175]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[175]) );
  d_ff \sig_prgm_register/genblk1[174].single_DFF  ( .d(
        \sig_prgm_register/or_signal [174]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[174]) );
  d_ff \sig_prgm_register/genblk1[173].single_DFF  ( .d(
        \sig_prgm_register/or_signal [173]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[173]) );
  d_ff \sig_prgm_register/genblk1[172].single_DFF  ( .d(
        \sig_prgm_register/or_signal [172]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[172]) );
  d_ff \sig_prgm_register/genblk1[171].single_DFF  ( .d(
        \sig_prgm_register/or_signal [171]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[171]) );
  d_ff \sig_prgm_register/genblk1[170].single_DFF  ( .d(
        \sig_prgm_register/or_signal [170]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[170]) );
  d_ff \sig_prgm_register/genblk1[169].single_DFF  ( .d(
        \sig_prgm_register/or_signal [169]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[169]) );
  d_ff \sig_prgm_register/genblk1[168].single_DFF  ( .d(
        \sig_prgm_register/or_signal [168]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[168]) );
  d_ff \sig_prgm_register/genblk1[167].single_DFF  ( .d(
        \sig_prgm_register/or_signal [167]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[167]) );
  d_ff \sig_prgm_register/genblk1[166].single_DFF  ( .d(
        \sig_prgm_register/or_signal [166]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[166]) );
  d_ff \sig_prgm_register/genblk1[165].single_DFF  ( .d(
        \sig_prgm_register/or_signal [165]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[165]) );
  d_ff \sig_prgm_register/genblk1[164].single_DFF  ( .d(
        \sig_prgm_register/or_signal [164]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[164]) );
  d_ff \sig_prgm_register/genblk1[163].single_DFF  ( .d(
        \sig_prgm_register/or_signal [163]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[163]) );
  d_ff \sig_prgm_register/genblk1[162].single_DFF  ( .d(
        \sig_prgm_register/or_signal [162]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[162]) );
  d_ff \sig_prgm_register/genblk1[161].single_DFF  ( .d(
        \sig_prgm_register/or_signal [161]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[161]) );
  d_ff \sig_prgm_register/genblk1[160].single_DFF  ( .d(
        \sig_prgm_register/or_signal [160]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[160]) );
  d_ff \sig_prgm_register/genblk1[159].single_DFF  ( .d(
        \sig_prgm_register/or_signal [159]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[159]) );
  d_ff \sig_prgm_register/genblk1[158].single_DFF  ( .d(
        \sig_prgm_register/or_signal [158]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[158]) );
  d_ff \sig_prgm_register/genblk1[157].single_DFF  ( .d(
        \sig_prgm_register/or_signal [157]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[157]) );
  d_ff \sig_prgm_register/genblk1[156].single_DFF  ( .d(
        \sig_prgm_register/or_signal [156]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[156]) );
  d_ff \sig_prgm_register/genblk1[155].single_DFF  ( .d(
        \sig_prgm_register/or_signal [155]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[155]) );
  d_ff \sig_prgm_register/genblk1[154].single_DFF  ( .d(
        \sig_prgm_register/or_signal [154]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[154]) );
  d_ff \sig_prgm_register/genblk1[153].single_DFF  ( .d(
        \sig_prgm_register/or_signal [153]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[153]) );
  d_ff \sig_prgm_register/genblk1[152].single_DFF  ( .d(
        \sig_prgm_register/or_signal [152]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[152]) );
  d_ff \sig_prgm_register/genblk1[151].single_DFF  ( .d(
        \sig_prgm_register/or_signal [151]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[151]) );
  d_ff \sig_prgm_register/genblk1[150].single_DFF  ( .d(
        \sig_prgm_register/or_signal [150]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[150]) );
  d_ff \sig_prgm_register/genblk1[149].single_DFF  ( .d(
        \sig_prgm_register/or_signal [149]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[149]) );
  d_ff \sig_prgm_register/genblk1[148].single_DFF  ( .d(
        \sig_prgm_register/or_signal [148]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[148]) );
  d_ff \sig_prgm_register/genblk1[147].single_DFF  ( .d(
        \sig_prgm_register/or_signal [147]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[147]) );
  d_ff \sig_prgm_register/genblk1[146].single_DFF  ( .d(
        \sig_prgm_register/or_signal [146]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[146]) );
  d_ff \sig_prgm_register/genblk1[145].single_DFF  ( .d(
        \sig_prgm_register/or_signal [145]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[145]) );
  d_ff \sig_prgm_register/genblk1[144].single_DFF  ( .d(
        \sig_prgm_register/or_signal [144]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[144]) );
  d_ff \sig_prgm_register/genblk1[143].single_DFF  ( .d(
        \sig_prgm_register/or_signal [143]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[143]) );
  d_ff \sig_prgm_register/genblk1[142].single_DFF  ( .d(
        \sig_prgm_register/or_signal [142]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[142]) );
  d_ff \sig_prgm_register/genblk1[141].single_DFF  ( .d(
        \sig_prgm_register/or_signal [141]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[141]) );
  d_ff \sig_prgm_register/genblk1[140].single_DFF  ( .d(
        \sig_prgm_register/or_signal [140]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[140]) );
  d_ff \sig_prgm_register/genblk1[139].single_DFF  ( .d(
        \sig_prgm_register/or_signal [139]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[139]) );
  d_ff \sig_prgm_register/genblk1[138].single_DFF  ( .d(
        \sig_prgm_register/or_signal [138]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[138]) );
  d_ff \sig_prgm_register/genblk1[137].single_DFF  ( .d(
        \sig_prgm_register/or_signal [137]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[137]) );
  d_ff \sig_prgm_register/genblk1[136].single_DFF  ( .d(
        \sig_prgm_register/or_signal [136]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[136]) );
  d_ff \sig_prgm_register/genblk1[135].single_DFF  ( .d(
        \sig_prgm_register/or_signal [135]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[135]) );
  d_ff \sig_prgm_register/genblk1[134].single_DFF  ( .d(
        \sig_prgm_register/or_signal [134]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[134]) );
  d_ff \sig_prgm_register/genblk1[133].single_DFF  ( .d(
        \sig_prgm_register/or_signal [133]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[133]) );
  d_ff \sig_prgm_register/genblk1[132].single_DFF  ( .d(
        \sig_prgm_register/or_signal [132]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[132]) );
  d_ff \sig_prgm_register/genblk1[131].single_DFF  ( .d(
        \sig_prgm_register/or_signal [131]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[131]) );
  d_ff \sig_prgm_register/genblk1[130].single_DFF  ( .d(
        \sig_prgm_register/or_signal [130]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[130]) );
  d_ff \sig_prgm_register/genblk1[129].single_DFF  ( .d(
        \sig_prgm_register/or_signal [129]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[129]) );
  d_ff \sig_prgm_register/genblk1[128].single_DFF  ( .d(
        \sig_prgm_register/or_signal [128]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[128]) );
  d_ff \sig_prgm_register/genblk1[127].single_DFF  ( .d(
        \sig_prgm_register/or_signal [127]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[127]) );
  d_ff \sig_prgm_register/genblk1[126].single_DFF  ( .d(
        \sig_prgm_register/or_signal [126]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[126]) );
  d_ff \sig_prgm_register/genblk1[125].single_DFF  ( .d(
        \sig_prgm_register/or_signal [125]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[125]) );
  d_ff \sig_prgm_register/genblk1[124].single_DFF  ( .d(
        \sig_prgm_register/or_signal [124]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[124]) );
  d_ff \sig_prgm_register/genblk1[123].single_DFF  ( .d(
        \sig_prgm_register/or_signal [123]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[123]) );
  d_ff \sig_prgm_register/genblk1[122].single_DFF  ( .d(
        \sig_prgm_register/or_signal [122]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[122]) );
  d_ff \sig_prgm_register/genblk1[121].single_DFF  ( .d(
        \sig_prgm_register/or_signal [121]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[121]) );
  d_ff \sig_prgm_register/genblk1[120].single_DFF  ( .d(
        \sig_prgm_register/or_signal [120]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[120]) );
  d_ff \sig_prgm_register/genblk1[119].single_DFF  ( .d(
        \sig_prgm_register/or_signal [119]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[119]) );
  d_ff \sig_prgm_register/genblk1[118].single_DFF  ( .d(
        \sig_prgm_register/or_signal [118]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[118]) );
  d_ff \sig_prgm_register/genblk1[117].single_DFF  ( .d(
        \sig_prgm_register/or_signal [117]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[117]) );
  d_ff \sig_prgm_register/genblk1[116].single_DFF  ( .d(
        \sig_prgm_register/or_signal [116]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[116]) );
  d_ff \sig_prgm_register/genblk1[115].single_DFF  ( .d(
        \sig_prgm_register/or_signal [115]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[115]) );
  d_ff \sig_prgm_register/genblk1[114].single_DFF  ( .d(
        \sig_prgm_register/or_signal [114]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[114]) );
  d_ff \sig_prgm_register/genblk1[113].single_DFF  ( .d(
        \sig_prgm_register/or_signal [113]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[113]) );
  d_ff \sig_prgm_register/genblk1[112].single_DFF  ( .d(
        \sig_prgm_register/or_signal [112]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[112]) );
  d_ff \sig_prgm_register/genblk1[111].single_DFF  ( .d(
        \sig_prgm_register/or_signal [111]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[111]) );
  d_ff \sig_prgm_register/genblk1[110].single_DFF  ( .d(
        \sig_prgm_register/or_signal [110]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[110]) );
  d_ff \sig_prgm_register/genblk1[109].single_DFF  ( .d(
        \sig_prgm_register/or_signal [109]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[109]) );
  d_ff \sig_prgm_register/genblk1[108].single_DFF  ( .d(
        \sig_prgm_register/or_signal [108]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[108]) );
  d_ff \sig_prgm_register/genblk1[107].single_DFF  ( .d(
        \sig_prgm_register/or_signal [107]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[107]) );
  d_ff \sig_prgm_register/genblk1[106].single_DFF  ( .d(
        \sig_prgm_register/or_signal [106]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[106]) );
  d_ff \sig_prgm_register/genblk1[105].single_DFF  ( .d(
        \sig_prgm_register/or_signal [105]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[105]) );
  d_ff \sig_prgm_register/genblk1[104].single_DFF  ( .d(
        \sig_prgm_register/or_signal [104]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[104]) );
  d_ff \sig_prgm_register/genblk1[103].single_DFF  ( .d(
        \sig_prgm_register/or_signal [103]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[103]) );
  d_ff \sig_prgm_register/genblk1[102].single_DFF  ( .d(
        \sig_prgm_register/or_signal [102]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[102]) );
  d_ff \sig_prgm_register/genblk1[101].single_DFF  ( .d(
        \sig_prgm_register/or_signal [101]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[101]) );
  d_ff \sig_prgm_register/genblk1[100].single_DFF  ( .d(
        \sig_prgm_register/or_signal [100]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[100]) );
  d_ff \sig_prgm_register/genblk1[99].single_DFF  ( .d(
        \sig_prgm_register/or_signal [99]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[99]) );
  d_ff \sig_prgm_register/genblk1[98].single_DFF  ( .d(
        \sig_prgm_register/or_signal [98]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[98]) );
  d_ff \sig_prgm_register/genblk1[97].single_DFF  ( .d(
        \sig_prgm_register/or_signal [97]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[97]) );
  d_ff \sig_prgm_register/genblk1[96].single_DFF  ( .d(
        \sig_prgm_register/or_signal [96]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[96]) );
  d_ff \sig_prgm_register/genblk1[95].single_DFF  ( .d(
        \sig_prgm_register/or_signal [95]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[95]) );
  d_ff \sig_prgm_register/genblk1[94].single_DFF  ( .d(
        \sig_prgm_register/or_signal [94]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[94]) );
  d_ff \sig_prgm_register/genblk1[93].single_DFF  ( .d(
        \sig_prgm_register/or_signal [93]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[93]) );
  d_ff \sig_prgm_register/genblk1[92].single_DFF  ( .d(
        \sig_prgm_register/or_signal [92]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[92]) );
  d_ff \sig_prgm_register/genblk1[91].single_DFF  ( .d(
        \sig_prgm_register/or_signal [91]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[91]) );
  d_ff \sig_prgm_register/genblk1[90].single_DFF  ( .d(
        \sig_prgm_register/or_signal [90]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[90]) );
  d_ff \sig_prgm_register/genblk1[89].single_DFF  ( .d(
        \sig_prgm_register/or_signal [89]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[89]) );
  d_ff \sig_prgm_register/genblk1[88].single_DFF  ( .d(
        \sig_prgm_register/or_signal [88]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[88]) );
  d_ff \sig_prgm_register/genblk1[87].single_DFF  ( .d(
        \sig_prgm_register/or_signal [87]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[87]) );
  d_ff \sig_prgm_register/genblk1[86].single_DFF  ( .d(
        \sig_prgm_register/or_signal [86]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[86]) );
  d_ff \sig_prgm_register/genblk1[85].single_DFF  ( .d(
        \sig_prgm_register/or_signal [85]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[85]) );
  d_ff \sig_prgm_register/genblk1[84].single_DFF  ( .d(
        \sig_prgm_register/or_signal [84]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[84]) );
  d_ff \sig_prgm_register/genblk1[83].single_DFF  ( .d(
        \sig_prgm_register/or_signal [83]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[83]) );
  d_ff \sig_prgm_register/genblk1[82].single_DFF  ( .d(
        \sig_prgm_register/or_signal [82]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[82]) );
  d_ff \sig_prgm_register/genblk1[81].single_DFF  ( .d(
        \sig_prgm_register/or_signal [81]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[81]) );
  d_ff \sig_prgm_register/genblk1[80].single_DFF  ( .d(
        \sig_prgm_register/or_signal [80]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[80]) );
  d_ff \sig_prgm_register/genblk1[79].single_DFF  ( .d(
        \sig_prgm_register/or_signal [79]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[79]) );
  d_ff \sig_prgm_register/genblk1[78].single_DFF  ( .d(
        \sig_prgm_register/or_signal [78]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[78]) );
  d_ff \sig_prgm_register/genblk1[77].single_DFF  ( .d(
        \sig_prgm_register/or_signal [77]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[77]) );
  d_ff \sig_prgm_register/genblk1[76].single_DFF  ( .d(
        \sig_prgm_register/or_signal [76]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[76]) );
  d_ff \sig_prgm_register/genblk1[75].single_DFF  ( .d(
        \sig_prgm_register/or_signal [75]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[75]) );
  d_ff \sig_prgm_register/genblk1[74].single_DFF  ( .d(
        \sig_prgm_register/or_signal [74]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[74]) );
  d_ff \sig_prgm_register/genblk1[73].single_DFF  ( .d(
        \sig_prgm_register/or_signal [73]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[73]) );
  d_ff \sig_prgm_register/genblk1[72].single_DFF  ( .d(
        \sig_prgm_register/or_signal [72]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[72]) );
  d_ff \sig_prgm_register/genblk1[71].single_DFF  ( .d(
        \sig_prgm_register/or_signal [71]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[71]) );
  d_ff \sig_prgm_register/genblk1[70].single_DFF  ( .d(
        \sig_prgm_register/or_signal [70]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[70]) );
  d_ff \sig_prgm_register/genblk1[69].single_DFF  ( .d(
        \sig_prgm_register/or_signal [69]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[69]) );
  d_ff \sig_prgm_register/genblk1[68].single_DFF  ( .d(
        \sig_prgm_register/or_signal [68]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[68]) );
  d_ff \sig_prgm_register/genblk1[67].single_DFF  ( .d(
        \sig_prgm_register/or_signal [67]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[67]) );
  d_ff \sig_prgm_register/genblk1[66].single_DFF  ( .d(
        \sig_prgm_register/or_signal [66]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[66]) );
  d_ff \sig_prgm_register/genblk1[65].single_DFF  ( .d(
        \sig_prgm_register/or_signal [65]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[65]) );
  d_ff \sig_prgm_register/genblk1[64].single_DFF  ( .d(
        \sig_prgm_register/or_signal [64]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[64]) );
  d_ff \sig_prgm_register/genblk1[63].single_DFF  ( .d(
        \sig_prgm_register/or_signal [63]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[63]) );
  d_ff \sig_prgm_register/genblk1[62].single_DFF  ( .d(
        \sig_prgm_register/or_signal [62]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[62]) );
  d_ff \sig_prgm_register/genblk1[61].single_DFF  ( .d(
        \sig_prgm_register/or_signal [61]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[61]) );
  d_ff \sig_prgm_register/genblk1[60].single_DFF  ( .d(
        \sig_prgm_register/or_signal [60]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[60]) );
  d_ff \sig_prgm_register/genblk1[59].single_DFF  ( .d(
        \sig_prgm_register/or_signal [59]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[59]) );
  d_ff \sig_prgm_register/genblk1[58].single_DFF  ( .d(
        \sig_prgm_register/or_signal [58]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[58]) );
  d_ff \sig_prgm_register/genblk1[57].single_DFF  ( .d(
        \sig_prgm_register/or_signal [57]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[57]) );
  d_ff \sig_prgm_register/genblk1[56].single_DFF  ( .d(
        \sig_prgm_register/or_signal [56]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[56]) );
  d_ff \sig_prgm_register/genblk1[55].single_DFF  ( .d(
        \sig_prgm_register/or_signal [55]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[55]) );
  d_ff \sig_prgm_register/genblk1[54].single_DFF  ( .d(
        \sig_prgm_register/or_signal [54]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[54]) );
  d_ff \sig_prgm_register/genblk1[53].single_DFF  ( .d(
        \sig_prgm_register/or_signal [53]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[53]) );
  d_ff \sig_prgm_register/genblk1[52].single_DFF  ( .d(
        \sig_prgm_register/or_signal [52]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[52]) );
  d_ff \sig_prgm_register/genblk1[51].single_DFF  ( .d(
        \sig_prgm_register/or_signal [51]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[51]) );
  d_ff \sig_prgm_register/genblk1[50].single_DFF  ( .d(
        \sig_prgm_register/or_signal [50]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[50]) );
  d_ff \sig_prgm_register/genblk1[49].single_DFF  ( .d(
        \sig_prgm_register/or_signal [49]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[49]) );
  d_ff \sig_prgm_register/genblk1[48].single_DFF  ( .d(
        \sig_prgm_register/or_signal [48]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[48]) );
  d_ff \sig_prgm_register/genblk1[47].single_DFF  ( .d(
        \sig_prgm_register/or_signal [47]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[47]) );
  d_ff \sig_prgm_register/genblk1[46].single_DFF  ( .d(
        \sig_prgm_register/or_signal [46]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[46]) );
  d_ff \sig_prgm_register/genblk1[45].single_DFF  ( .d(
        \sig_prgm_register/or_signal [45]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[45]) );
  d_ff \sig_prgm_register/genblk1[44].single_DFF  ( .d(
        \sig_prgm_register/or_signal [44]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[44]) );
  d_ff \sig_prgm_register/genblk1[43].single_DFF  ( .d(
        \sig_prgm_register/or_signal [43]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[43]) );
  d_ff \sig_prgm_register/genblk1[42].single_DFF  ( .d(
        \sig_prgm_register/or_signal [42]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[42]) );
  d_ff \sig_prgm_register/genblk1[41].single_DFF  ( .d(
        \sig_prgm_register/or_signal [41]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[41]) );
  d_ff \sig_prgm_register/genblk1[40].single_DFF  ( .d(
        \sig_prgm_register/or_signal [40]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[40]) );
  d_ff \sig_prgm_register/genblk1[39].single_DFF  ( .d(
        \sig_prgm_register/or_signal [39]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[39]) );
  d_ff \sig_prgm_register/genblk1[38].single_DFF  ( .d(
        \sig_prgm_register/or_signal [38]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[38]) );
  d_ff \sig_prgm_register/genblk1[37].single_DFF  ( .d(
        \sig_prgm_register/or_signal [37]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[37]) );
  d_ff \sig_prgm_register/genblk1[36].single_DFF  ( .d(
        \sig_prgm_register/or_signal [36]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[36]) );
  d_ff \sig_prgm_register/genblk1[35].single_DFF  ( .d(
        \sig_prgm_register/or_signal [35]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[35]) );
  d_ff \sig_prgm_register/genblk1[34].single_DFF  ( .d(
        \sig_prgm_register/or_signal [34]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[34]) );
  d_ff \sig_prgm_register/genblk1[33].single_DFF  ( .d(
        \sig_prgm_register/or_signal [33]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[33]) );
  d_ff \sig_prgm_register/genblk1[32].single_DFF  ( .d(
        \sig_prgm_register/or_signal [32]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[32]) );
  d_ff \sig_prgm_register/genblk1[31].single_DFF  ( .d(
        \sig_prgm_register/or_signal [31]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[31]) );
  d_ff \sig_prgm_register/genblk1[30].single_DFF  ( .d(
        \sig_prgm_register/or_signal [30]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[30]) );
  d_ff \sig_prgm_register/genblk1[29].single_DFF  ( .d(
        \sig_prgm_register/or_signal [29]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[29]) );
  d_ff \sig_prgm_register/genblk1[28].single_DFF  ( .d(
        \sig_prgm_register/or_signal [28]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[28]) );
  d_ff \sig_prgm_register/genblk1[27].single_DFF  ( .d(
        \sig_prgm_register/or_signal [27]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[27]) );
  d_ff \sig_prgm_register/genblk1[26].single_DFF  ( .d(
        \sig_prgm_register/or_signal [26]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[26]) );
  d_ff \sig_prgm_register/genblk1[25].single_DFF  ( .d(
        \sig_prgm_register/or_signal [25]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[25]) );
  d_ff \sig_prgm_register/genblk1[24].single_DFF  ( .d(
        \sig_prgm_register/or_signal [24]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[24]) );
  d_ff \sig_prgm_register/genblk1[23].single_DFF  ( .d(
        \sig_prgm_register/or_signal [23]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[23]) );
  d_ff \sig_prgm_register/genblk1[22].single_DFF  ( .d(
        \sig_prgm_register/or_signal [22]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[22]) );
  d_ff \sig_prgm_register/genblk1[21].single_DFF  ( .d(
        \sig_prgm_register/or_signal [21]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[21]) );
  d_ff \sig_prgm_register/genblk1[20].single_DFF  ( .d(
        \sig_prgm_register/or_signal [20]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[20]) );
  d_ff \sig_prgm_register/genblk1[19].single_DFF  ( .d(
        \sig_prgm_register/or_signal [19]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[19]) );
  d_ff \sig_prgm_register/genblk1[18].single_DFF  ( .d(
        \sig_prgm_register/or_signal [18]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[18]) );
  d_ff \sig_prgm_register/genblk1[17].single_DFF  ( .d(
        \sig_prgm_register/or_signal [17]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[17]) );
  d_ff \sig_prgm_register/genblk1[16].single_DFF  ( .d(
        \sig_prgm_register/or_signal [16]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[16]) );
  d_ff \sig_prgm_register/genblk1[15].single_DFF  ( .d(
        \sig_prgm_register/or_signal [15]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[15]) );
  d_ff \sig_prgm_register/genblk1[14].single_DFF  ( .d(
        \sig_prgm_register/or_signal [14]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[14]) );
  d_ff \sig_prgm_register/genblk1[13].single_DFF  ( .d(
        \sig_prgm_register/or_signal [13]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[13]) );
  d_ff \sig_prgm_register/genblk1[12].single_DFF  ( .d(
        \sig_prgm_register/or_signal [12]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[12]) );
  d_ff \sig_prgm_register/genblk1[11].single_DFF  ( .d(
        \sig_prgm_register/or_signal [11]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[11]) );
  d_ff \sig_prgm_register/genblk1[10].single_DFF  ( .d(
        \sig_prgm_register/or_signal [10]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[10]) );
  d_ff \sig_prgm_register/genblk1[9].single_DFF  ( .d(
        \sig_prgm_register/or_signal [9]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[9]) );
  d_ff \sig_prgm_register/genblk1[8].single_DFF  ( .d(
        \sig_prgm_register/or_signal [8]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[8]) );
  d_ff \sig_prgm_register/genblk1[7].single_DFF  ( .d(
        \sig_prgm_register/or_signal [7]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[7]) );
  d_ff \sig_prgm_register/genblk1[6].single_DFF  ( .d(
        \sig_prgm_register/or_signal [6]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[6]) );
  d_ff \sig_prgm_register/genblk1[5].single_DFF  ( .d(
        \sig_prgm_register/or_signal [5]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[5]) );
  d_ff \sig_prgm_register/genblk1[4].single_DFF  ( .d(
        \sig_prgm_register/or_signal [4]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[4]) );
  d_ff \sig_prgm_register/genblk1[3].single_DFF  ( .d(
        \sig_prgm_register/or_signal [3]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[3]) );
  d_ff \sig_prgm_register/genblk1[2].single_DFF  ( .d(
        \sig_prgm_register/or_signal [2]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[2]) );
  d_ff \sig_prgm_register/genblk1[1].single_DFF  ( .d(
        \sig_prgm_register/or_signal [1]), .clk(clk), .R(
        \sig_prgm_register/clear_not ), .Q(b[1]) );
  d_ff \sig_prgm_register/first_DFF  ( .d(\sig_prgm_register/or_signal [0]), 
        .clk(clk), .R(\sig_prgm_register/clear_not ), .Q(b[0]) );
  inv U2 ( .a(n1), .out(\sig_prgm_register/or_signal [0]) );
  inv U3 ( .a(n2), .out(\sig_prgm_register/or_signal [1]) );
  inv U4 ( .a(n3), .out(\sig_prgm_register/or_signal [2]) );
  inv U5 ( .a(n4), .out(\sig_prgm_register/or_signal [3]) );
  inv U6 ( .a(n5), .out(\sig_prgm_register/or_signal [4]) );
  inv U7 ( .a(n6), .out(\sig_prgm_register/or_signal [5]) );
  inv U8 ( .a(n7), .out(\sig_prgm_register/or_signal [6]) );
  inv U9 ( .a(n8), .out(\sig_prgm_register/or_signal [7]) );
  inv U10 ( .a(n9), .out(\sig_prgm_register/or_signal [8]) );
  inv U11 ( .a(n10), .out(\sig_prgm_register/or_signal [9]) );
  inv U12 ( .a(n11), .out(\sig_prgm_register/or_signal [10]) );
  inv U13 ( .a(n12), .out(\sig_prgm_register/or_signal [11]) );
  inv U14 ( .a(n13), .out(\sig_prgm_register/or_signal [12]) );
  inv U15 ( .a(n14), .out(\sig_prgm_register/or_signal [13]) );
  inv U16 ( .a(n15), .out(\sig_prgm_register/or_signal [14]) );
  inv U17 ( .a(n16), .out(\sig_prgm_register/or_signal [15]) );
  inv U18 ( .a(n17), .out(\sig_prgm_register/or_signal [16]) );
  inv U19 ( .a(n18), .out(\sig_prgm_register/or_signal [17]) );
  inv U20 ( .a(n19), .out(\sig_prgm_register/or_signal [18]) );
  inv U21 ( .a(n20), .out(\sig_prgm_register/or_signal [19]) );
  inv U22 ( .a(n21), .out(\sig_prgm_register/or_signal [20]) );
  inv U23 ( .a(n22), .out(\sig_prgm_register/or_signal [21]) );
  inv U24 ( .a(n23), .out(\sig_prgm_register/or_signal [22]) );
  inv U25 ( .a(n24), .out(\sig_prgm_register/or_signal [23]) );
  inv U26 ( .a(n25), .out(\sig_prgm_register/or_signal [24]) );
  inv U27 ( .a(n26), .out(\sig_prgm_register/or_signal [25]) );
  inv U28 ( .a(n27), .out(\sig_prgm_register/or_signal [26]) );
  inv U29 ( .a(n28), .out(\sig_prgm_register/or_signal [27]) );
  inv U30 ( .a(n29), .out(\sig_prgm_register/or_signal [28]) );
  inv U31 ( .a(n30), .out(\sig_prgm_register/or_signal [29]) );
  inv U32 ( .a(n31), .out(\sig_prgm_register/or_signal [30]) );
  inv U33 ( .a(n32), .out(\sig_prgm_register/or_signal [31]) );
  inv U34 ( .a(n33), .out(\sig_prgm_register/or_signal [32]) );
  inv U35 ( .a(n34), .out(\sig_prgm_register/or_signal [33]) );
  inv U36 ( .a(n35), .out(\sig_prgm_register/or_signal [34]) );
  inv U37 ( .a(n36), .out(\sig_prgm_register/or_signal [35]) );
  inv U38 ( .a(n37), .out(\sig_prgm_register/or_signal [36]) );
  inv U39 ( .a(n38), .out(\sig_prgm_register/or_signal [37]) );
  inv U40 ( .a(n39), .out(\sig_prgm_register/or_signal [38]) );
  inv U41 ( .a(n40), .out(\sig_prgm_register/or_signal [39]) );
  inv U42 ( .a(n41), .out(\sig_prgm_register/or_signal [40]) );
  inv U43 ( .a(n42), .out(\sig_prgm_register/or_signal [41]) );
  inv U44 ( .a(n43), .out(\sig_prgm_register/or_signal [42]) );
  inv U45 ( .a(n44), .out(\sig_prgm_register/or_signal [43]) );
  inv U46 ( .a(n45), .out(\sig_prgm_register/or_signal [44]) );
  inv U47 ( .a(n46), .out(\sig_prgm_register/or_signal [45]) );
  inv U48 ( .a(n47), .out(\sig_prgm_register/or_signal [46]) );
  inv U49 ( .a(n48), .out(\sig_prgm_register/or_signal [47]) );
  inv U50 ( .a(n49), .out(\sig_prgm_register/or_signal [48]) );
  inv U51 ( .a(n50), .out(\sig_prgm_register/or_signal [49]) );
  inv U52 ( .a(n51), .out(\sig_prgm_register/or_signal [50]) );
  inv U53 ( .a(n52), .out(\sig_prgm_register/or_signal [51]) );
  inv U54 ( .a(n53), .out(\sig_prgm_register/or_signal [52]) );
  inv U55 ( .a(n54), .out(\sig_prgm_register/or_signal [53]) );
  inv U56 ( .a(n55), .out(\sig_prgm_register/or_signal [54]) );
  inv U57 ( .a(n56), .out(\sig_prgm_register/or_signal [55]) );
  inv U58 ( .a(n57), .out(\sig_prgm_register/or_signal [56]) );
  inv U59 ( .a(n58), .out(\sig_prgm_register/or_signal [57]) );
  inv U60 ( .a(n59), .out(\sig_prgm_register/or_signal [58]) );
  inv U61 ( .a(n60), .out(\sig_prgm_register/or_signal [59]) );
  inv U62 ( .a(n61), .out(\sig_prgm_register/or_signal [60]) );
  inv U63 ( .a(n62), .out(\sig_prgm_register/or_signal [61]) );
  inv U64 ( .a(n63), .out(\sig_prgm_register/or_signal [62]) );
  inv U65 ( .a(n64), .out(\sig_prgm_register/or_signal [63]) );
  inv U66 ( .a(n65), .out(\sig_prgm_register/or_signal [64]) );
  inv U67 ( .a(n66), .out(\sig_prgm_register/or_signal [65]) );
  inv U68 ( .a(n67), .out(\sig_prgm_register/or_signal [66]) );
  inv U69 ( .a(n68), .out(\sig_prgm_register/or_signal [67]) );
  inv U70 ( .a(n69), .out(\sig_prgm_register/or_signal [68]) );
  inv U71 ( .a(n70), .out(\sig_prgm_register/or_signal [69]) );
  inv U72 ( .a(n71), .out(\sig_prgm_register/or_signal [70]) );
  inv U73 ( .a(n72), .out(\sig_prgm_register/or_signal [71]) );
  inv U74 ( .a(n73), .out(\sig_prgm_register/or_signal [72]) );
  inv U75 ( .a(n74), .out(\sig_prgm_register/or_signal [73]) );
  inv U76 ( .a(n75), .out(\sig_prgm_register/or_signal [74]) );
  inv U77 ( .a(n76), .out(\sig_prgm_register/or_signal [75]) );
  inv U78 ( .a(n77), .out(\sig_prgm_register/or_signal [76]) );
  inv U79 ( .a(n78), .out(\sig_prgm_register/or_signal [77]) );
  inv U80 ( .a(n79), .out(\sig_prgm_register/or_signal [78]) );
  inv U81 ( .a(n80), .out(\sig_prgm_register/or_signal [79]) );
  inv U82 ( .a(n81), .out(\sig_prgm_register/or_signal [80]) );
  inv U83 ( .a(n82), .out(\sig_prgm_register/or_signal [81]) );
  inv U84 ( .a(n83), .out(\sig_prgm_register/or_signal [82]) );
  inv U85 ( .a(n84), .out(\sig_prgm_register/or_signal [83]) );
  inv U86 ( .a(n85), .out(\sig_prgm_register/or_signal [84]) );
  inv U87 ( .a(n86), .out(\sig_prgm_register/or_signal [85]) );
  inv U88 ( .a(n87), .out(\sig_prgm_register/or_signal [86]) );
  inv U89 ( .a(n88), .out(\sig_prgm_register/or_signal [87]) );
  inv U90 ( .a(n89), .out(\sig_prgm_register/or_signal [88]) );
  inv U91 ( .a(n90), .out(\sig_prgm_register/or_signal [89]) );
  inv U92 ( .a(n91), .out(\sig_prgm_register/or_signal [90]) );
  inv U93 ( .a(n92), .out(\sig_prgm_register/or_signal [91]) );
  inv U94 ( .a(n93), .out(\sig_prgm_register/or_signal [92]) );
  inv U95 ( .a(n94), .out(\sig_prgm_register/or_signal [93]) );
  inv U96 ( .a(n95), .out(\sig_prgm_register/or_signal [94]) );
  inv U97 ( .a(n96), .out(\sig_prgm_register/or_signal [95]) );
  inv U98 ( .a(n97), .out(\sig_prgm_register/or_signal [96]) );
  inv U99 ( .a(n98), .out(\sig_prgm_register/or_signal [97]) );
  inv U100 ( .a(n99), .out(\sig_prgm_register/or_signal [98]) );
  inv U101 ( .a(n100), .out(\sig_prgm_register/or_signal [99]) );
  inv U102 ( .a(n101), .out(\sig_prgm_register/or_signal [100]) );
  inv U103 ( .a(n102), .out(\sig_prgm_register/or_signal [101]) );
  inv U104 ( .a(n103), .out(\sig_prgm_register/or_signal [102]) );
  inv U105 ( .a(n104), .out(\sig_prgm_register/or_signal [103]) );
  inv U106 ( .a(n105), .out(\sig_prgm_register/or_signal [104]) );
  inv U107 ( .a(n106), .out(\sig_prgm_register/or_signal [105]) );
  inv U108 ( .a(n107), .out(\sig_prgm_register/or_signal [106]) );
  inv U109 ( .a(n108), .out(\sig_prgm_register/or_signal [107]) );
  inv U110 ( .a(n109), .out(\sig_prgm_register/or_signal [108]) );
  inv U111 ( .a(n110), .out(\sig_prgm_register/or_signal [109]) );
  inv U112 ( .a(n111), .out(\sig_prgm_register/or_signal [110]) );
  inv U113 ( .a(n112), .out(\sig_prgm_register/or_signal [111]) );
  inv U114 ( .a(n113), .out(\sig_prgm_register/or_signal [112]) );
  inv U115 ( .a(n114), .out(\sig_prgm_register/or_signal [113]) );
  inv U116 ( .a(n115), .out(\sig_prgm_register/or_signal [114]) );
  inv U117 ( .a(n116), .out(\sig_prgm_register/or_signal [115]) );
  inv U118 ( .a(n117), .out(\sig_prgm_register/or_signal [116]) );
  inv U119 ( .a(n118), .out(\sig_prgm_register/or_signal [117]) );
  inv U120 ( .a(n119), .out(\sig_prgm_register/or_signal [118]) );
  inv U121 ( .a(n120), .out(\sig_prgm_register/or_signal [119]) );
  inv U122 ( .a(n121), .out(\sig_prgm_register/or_signal [120]) );
  inv U123 ( .a(n122), .out(\sig_prgm_register/or_signal [121]) );
  inv U124 ( .a(n123), .out(\sig_prgm_register/or_signal [122]) );
  inv U125 ( .a(n124), .out(\sig_prgm_register/or_signal [123]) );
  inv U126 ( .a(n125), .out(\sig_prgm_register/or_signal [124]) );
  inv U127 ( .a(n126), .out(\sig_prgm_register/or_signal [125]) );
  inv U128 ( .a(n127), .out(\sig_prgm_register/or_signal [126]) );
  inv U129 ( .a(n128), .out(\sig_prgm_register/or_signal [127]) );
  inv U130 ( .a(n129), .out(\sig_prgm_register/or_signal [128]) );
  inv U131 ( .a(n130), .out(\sig_prgm_register/or_signal [129]) );
  inv U132 ( .a(n131), .out(\sig_prgm_register/or_signal [130]) );
  inv U133 ( .a(n132), .out(\sig_prgm_register/or_signal [131]) );
  inv U134 ( .a(n133), .out(\sig_prgm_register/or_signal [132]) );
  inv U135 ( .a(n134), .out(\sig_prgm_register/or_signal [133]) );
  inv U136 ( .a(n135), .out(\sig_prgm_register/or_signal [134]) );
  inv U137 ( .a(n136), .out(\sig_prgm_register/or_signal [135]) );
  inv U138 ( .a(n137), .out(\sig_prgm_register/or_signal [136]) );
  inv U139 ( .a(n138), .out(\sig_prgm_register/or_signal [137]) );
  inv U140 ( .a(n139), .out(\sig_prgm_register/or_signal [138]) );
  inv U141 ( .a(n140), .out(\sig_prgm_register/or_signal [139]) );
  inv U142 ( .a(n141), .out(\sig_prgm_register/or_signal [140]) );
  inv U143 ( .a(n142), .out(\sig_prgm_register/or_signal [141]) );
  inv U144 ( .a(n143), .out(\sig_prgm_register/or_signal [142]) );
  inv U145 ( .a(n144), .out(\sig_prgm_register/or_signal [143]) );
  inv U146 ( .a(n145), .out(\sig_prgm_register/or_signal [144]) );
  inv U147 ( .a(n146), .out(\sig_prgm_register/or_signal [145]) );
  inv U148 ( .a(n147), .out(\sig_prgm_register/or_signal [146]) );
  inv U149 ( .a(n148), .out(\sig_prgm_register/or_signal [147]) );
  inv U150 ( .a(n149), .out(\sig_prgm_register/or_signal [148]) );
  inv U151 ( .a(n150), .out(\sig_prgm_register/or_signal [149]) );
  inv U152 ( .a(n151), .out(\sig_prgm_register/or_signal [150]) );
  inv U153 ( .a(n152), .out(\sig_prgm_register/or_signal [151]) );
  inv U154 ( .a(n153), .out(\sig_prgm_register/or_signal [152]) );
  inv U155 ( .a(n154), .out(\sig_prgm_register/or_signal [153]) );
  inv U156 ( .a(n155), .out(\sig_prgm_register/or_signal [154]) );
  inv U157 ( .a(n156), .out(\sig_prgm_register/or_signal [155]) );
  inv U158 ( .a(n157), .out(\sig_prgm_register/or_signal [156]) );
  inv U159 ( .a(n158), .out(\sig_prgm_register/or_signal [157]) );
  inv U160 ( .a(n159), .out(\sig_prgm_register/or_signal [158]) );
  inv U161 ( .a(n160), .out(\sig_prgm_register/or_signal [159]) );
  inv U162 ( .a(n161), .out(\sig_prgm_register/or_signal [160]) );
  inv U163 ( .a(n162), .out(\sig_prgm_register/or_signal [161]) );
  inv U164 ( .a(n163), .out(\sig_prgm_register/or_signal [162]) );
  inv U165 ( .a(n164), .out(\sig_prgm_register/or_signal [163]) );
  inv U166 ( .a(n165), .out(\sig_prgm_register/or_signal [164]) );
  inv U167 ( .a(n166), .out(\sig_prgm_register/or_signal [165]) );
  inv U168 ( .a(n167), .out(\sig_prgm_register/or_signal [166]) );
  inv U169 ( .a(n168), .out(\sig_prgm_register/or_signal [167]) );
  inv U170 ( .a(n169), .out(\sig_prgm_register/or_signal [168]) );
  inv U171 ( .a(n170), .out(\sig_prgm_register/or_signal [169]) );
  inv U172 ( .a(n171), .out(\sig_prgm_register/or_signal [170]) );
  inv U173 ( .a(n172), .out(\sig_prgm_register/or_signal [171]) );
  inv U174 ( .a(n173), .out(\sig_prgm_register/or_signal [172]) );
  inv U175 ( .a(n174), .out(\sig_prgm_register/or_signal [173]) );
  inv U176 ( .a(n175), .out(\sig_prgm_register/or_signal [174]) );
  inv U177 ( .a(n176), .out(\sig_prgm_register/or_signal [175]) );
  inv U178 ( .a(n177), .out(\sig_prgm_register/or_signal [176]) );
  inv U179 ( .a(n178), .out(\sig_prgm_register/or_signal [177]) );
  inv U180 ( .a(n179), .out(\sig_prgm_register/or_signal [178]) );
  inv U181 ( .a(n180), .out(\sig_prgm_register/or_signal [179]) );
  inv U182 ( .a(n181), .out(\sig_prgm_register/or_signal [180]) );
  inv U183 ( .a(n182), .out(\sig_prgm_register/or_signal [181]) );
  inv U184 ( .a(n183), .out(\sig_prgm_register/or_signal [182]) );
  inv U185 ( .a(n184), .out(\sig_prgm_register/or_signal [183]) );
  inv U186 ( .a(n185), .out(\sig_prgm_register/or_signal [184]) );
  inv U187 ( .a(n186), .out(\sig_prgm_register/or_signal [185]) );
  inv U188 ( .a(n187), .out(\sig_prgm_register/or_signal [186]) );
  inv U189 ( .a(n188), .out(\sig_prgm_register/or_signal [187]) );
  inv U190 ( .a(n189), .out(\sig_prgm_register/or_signal [188]) );
  inv U191 ( .a(n190), .out(\sig_prgm_register/or_signal [189]) );
  inv U192 ( .a(n191), .out(\sig_prgm_register/or_signal [190]) );
  inv U193 ( .a(n192), .out(\sig_prgm_register/or_signal [191]) );
  inv U194 ( .a(n193), .out(\sig_prgm_register/or_signal [192]) );
  inv U195 ( .a(n194), .out(\sig_prgm_register/or_signal [193]) );
  inv U196 ( .a(n195), .out(\sig_prgm_register/or_signal [194]) );
  inv U197 ( .a(n196), .out(\sig_prgm_register/or_signal [195]) );
  inv U198 ( .a(n197), .out(\sig_prgm_register/or_signal [196]) );
  inv U199 ( .a(n198), .out(\sig_prgm_register/or_signal [197]) );
  inv U200 ( .a(n199), .out(\sig_prgm_register/or_signal [198]) );
  inv U201 ( .a(n200), .out(\sig_prgm_register/or_signal [199]) );
  inv U202 ( .a(n201), .out(\sig_prgm_register/or_signal [200]) );
  inv U203 ( .a(n202), .out(\sig_prgm_register/or_signal [201]) );
  inv U204 ( .a(n203), .out(\sig_prgm_register/or_signal [202]) );
  inv U205 ( .a(n204), .out(\sig_prgm_register/or_signal [203]) );
  inv U206 ( .a(n205), .out(\sig_prgm_register/or_signal [204]) );
  inv U207 ( .a(n206), .out(\sig_prgm_register/or_signal [205]) );
  inv U208 ( .a(n207), .out(\sig_prgm_register/or_signal [206]) );
  inv U209 ( .a(n208), .out(\sig_prgm_register/or_signal [207]) );
  inv U210 ( .a(n209), .out(\sig_prgm_register/or_signal [208]) );
  inv U211 ( .a(n210), .out(\sig_prgm_register/or_signal [209]) );
  inv U212 ( .a(n211), .out(\sig_prgm_register/or_signal [210]) );
  inv U213 ( .a(n212), .out(\sig_prgm_register/or_signal [211]) );
  inv U214 ( .a(n213), .out(\sig_prgm_register/or_signal [212]) );
  inv U215 ( .a(n214), .out(\sig_prgm_register/or_signal [213]) );
  inv U216 ( .a(n215), .out(\sig_prgm_register/or_signal [214]) );
  inv U217 ( .a(n216), .out(\sig_prgm_register/or_signal [215]) );
  inv U218 ( .a(n217), .out(\sig_prgm_register/or_signal [216]) );
  inv U219 ( .a(n218), .out(\sig_prgm_register/or_signal [217]) );
  inv U220 ( .a(n219), .out(\sig_prgm_register/or_signal [218]) );
  inv U221 ( .a(n220), .out(\sig_prgm_register/or_signal [219]) );
  inv U222 ( .a(n221), .out(\sig_prgm_register/or_signal [220]) );
  inv U223 ( .a(n222), .out(\sig_prgm_register/or_signal [221]) );
  inv U224 ( .a(n223), .out(\sig_prgm_register/or_signal [222]) );
  inv U225 ( .a(n224), .out(\sig_prgm_register/or_signal [223]) );
  inv U226 ( .a(n225), .out(\sig_prgm_register/or_signal [224]) );
  inv U227 ( .a(n226), .out(\sig_prgm_register/or_signal [225]) );
  inv U228 ( .a(n227), .out(\sig_prgm_register/or_signal [226]) );
  inv U229 ( .a(n228), .out(\sig_prgm_register/or_signal [227]) );
  inv U230 ( .a(n229), .out(\sig_prgm_register/or_signal [228]) );
  inv U231 ( .a(n230), .out(\sig_prgm_register/or_signal [229]) );
  inv U232 ( .a(n231), .out(\sig_prgm_register/or_signal [230]) );
  inv U233 ( .a(n232), .out(\sig_prgm_register/or_signal [231]) );
  inv U234 ( .a(n233), .out(\sig_prgm_register/or_signal [232]) );
  inv U235 ( .a(n234), .out(\sig_prgm_register/or_signal [233]) );
  inv U236 ( .a(n235), .out(\sig_prgm_register/or_signal [234]) );
  inv U237 ( .a(n236), .out(\sig_prgm_register/or_signal [235]) );
  inv U238 ( .a(n237), .out(\sig_prgm_register/or_signal [236]) );
  inv U239 ( .a(n238), .out(\sig_prgm_register/or_signal [237]) );
  inv U240 ( .a(n239), .out(\sig_prgm_register/or_signal [238]) );
  inv U241 ( .a(n240), .out(\sig_prgm_register/or_signal [239]) );
  inv U242 ( .a(n241), .out(\sig_prgm_register/or_signal [240]) );
  inv U243 ( .a(n242), .out(\sig_prgm_register/or_signal [241]) );
  inv U244 ( .a(n243), .out(\sig_prgm_register/or_signal [242]) );
  inv U245 ( .a(n244), .out(\sig_prgm_register/or_signal [243]) );
  inv U246 ( .a(n245), .out(\sig_prgm_register/or_signal [244]) );
  inv U247 ( .a(n246), .out(\sig_prgm_register/or_signal [245]) );
  inv U248 ( .a(n247), .out(\sig_prgm_register/or_signal [246]) );
  inv U249 ( .a(n248), .out(\sig_prgm_register/or_signal [247]) );
  inv U250 ( .a(n249), .out(\sig_prgm_register/or_signal [248]) );
  inv U251 ( .a(n250), .out(\sig_prgm_register/or_signal [249]) );
  inv U252 ( .a(n251), .out(\sig_prgm_register/or_signal [250]) );
  inv U253 ( .a(n252), .out(\sig_prgm_register/or_signal [251]) );
  inv U254 ( .a(n253), .out(\sig_prgm_register/or_signal [252]) );
  inv U255 ( .a(n254), .out(\sig_prgm_register/or_signal [253]) );
  inv U256 ( .a(n255), .out(\sig_prgm_register/or_signal [254]) );
  inv U257 ( .a(n256), .out(\sig_prgm_register/or_signal [255]) );
  inv U258 ( .a(n257), .out(\sig_prgm_register/or_signal [256]) );
  inv U259 ( .a(n258), .out(\sig_prgm_register/or_signal [257]) );
  inv U260 ( .a(n259), .out(\sig_prgm_register/or_signal [258]) );
  inv U261 ( .a(n260), .out(\sig_prgm_register/or_signal [259]) );
  inv U262 ( .a(n261), .out(\sig_prgm_register/or_signal [260]) );
  inv U263 ( .a(n262), .out(\sig_prgm_register/or_signal [261]) );
  inv U264 ( .a(n263), .out(\sig_prgm_register/or_signal [262]) );
  inv U265 ( .a(n264), .out(\sig_prgm_register/or_signal [263]) );
  inv U266 ( .a(n265), .out(\sig_prgm_register/or_signal [264]) );
  inv U267 ( .a(n266), .out(\sig_prgm_register/or_signal [265]) );
  inv U268 ( .a(n267), .out(\sig_prgm_register/or_signal [266]) );
  inv U269 ( .a(n268), .out(\sig_prgm_register/or_signal [267]) );
  inv U270 ( .a(n269), .out(\sig_prgm_register/or_signal [268]) );
  inv U271 ( .a(n270), .out(\sig_prgm_register/or_signal [269]) );
  inv U272 ( .a(n271), .out(\sig_prgm_register/or_signal [270]) );
  inv U273 ( .a(n272), .out(\sig_prgm_register/or_signal [271]) );
  inv U274 ( .a(n273), .out(\sig_prgm_register/or_signal [272]) );
  inv U275 ( .a(n274), .out(\sig_prgm_register/or_signal [273]) );
  inv U276 ( .a(n275), .out(\sig_prgm_register/or_signal [274]) );
  inv U277 ( .a(n276), .out(\sig_prgm_register/or_signal [275]) );
  inv U278 ( .a(n277), .out(\sig_prgm_register/or_signal [276]) );
  inv U279 ( .a(n278), .out(\sig_prgm_register/or_signal [277]) );
  inv U280 ( .a(n279), .out(\sig_prgm_register/or_signal [278]) );
  inv U281 ( .a(n280), .out(\sig_prgm_register/or_signal [279]) );
  inv U282 ( .a(n281), .out(\sig_prgm_register/or_signal [280]) );
  inv U283 ( .a(n282), .out(\sig_prgm_register/or_signal [281]) );
  inv U284 ( .a(n283), .out(\sig_prgm_register/or_signal [282]) );
  inv U285 ( .a(n284), .out(\sig_prgm_register/or_signal [283]) );
  inv U286 ( .a(n285), .out(\sig_prgm_register/or_signal [284]) );
  inv U287 ( .a(n286), .out(\sig_prgm_register/or_signal [285]) );
  inv U288 ( .a(n287), .out(\sig_prgm_register/or_signal [286]) );
  inv U289 ( .a(n288), .out(\sig_prgm_register/or_signal [287]) );
  inv U290 ( .a(n289), .out(\sig_prgm_register/or_signal [288]) );
  inv U291 ( .a(n290), .out(\sig_prgm_register/or_signal [289]) );
  inv U292 ( .a(n291), .out(\sig_prgm_register/or_signal [290]) );
  inv U293 ( .a(n292), .out(\sig_prgm_register/or_signal [291]) );
  inv U294 ( .a(n293), .out(\sig_prgm_register/or_signal [292]) );
  inv U295 ( .a(n294), .out(\sig_prgm_register/or_signal [293]) );
  inv U296 ( .a(n295), .out(\sig_prgm_register/or_signal [294]) );
  inv U297 ( .a(n296), .out(\sig_prgm_register/or_signal [295]) );
  inv U298 ( .a(n297), .out(\sig_prgm_register/or_signal [296]) );
  inv U299 ( .a(n298), .out(\sig_prgm_register/or_signal [297]) );
  inv U300 ( .a(n299), .out(\sig_prgm_register/or_signal [298]) );
  inv U301 ( .a(n300), .out(\sig_prgm_register/or_signal [299]) );
  inv U302 ( .a(n301), .out(\sig_prgm_register/or_signal [300]) );
  inv U303 ( .a(n302), .out(\sig_prgm_register/or_signal [301]) );
  inv U304 ( .a(n303), .out(\sig_prgm_register/or_signal [302]) );
  inv U305 ( .a(n304), .out(\sig_prgm_register/or_signal [303]) );
  inv U306 ( .a(n305), .out(\sig_prgm_register/or_signal [304]) );
  inv U307 ( .a(n306), .out(\sig_prgm_register/or_signal [305]) );
  inv U308 ( .a(n307), .out(\sig_prgm_register/or_signal [306]) );
  inv U309 ( .a(n308), .out(\sig_prgm_register/or_signal [307]) );
  inv U310 ( .a(n309), .out(\sig_prgm_register/or_signal [308]) );
  inv U311 ( .a(n310), .out(\sig_prgm_register/or_signal [309]) );
  inv U312 ( .a(n311), .out(\sig_prgm_register/or_signal [310]) );
  inv U313 ( .a(n312), .out(\sig_prgm_register/or_signal [311]) );
  inv U314 ( .a(n313), .out(\sig_prgm_register/or_signal [312]) );
  inv U315 ( .a(n314), .out(\sig_prgm_register/or_signal [313]) );
  inv U316 ( .a(n315), .out(\sig_prgm_register/or_signal [314]) );
  inv U317 ( .a(n316), .out(\sig_prgm_register/or_signal [315]) );
  inv U318 ( .a(n317), .out(\sig_prgm_register/or_signal [316]) );
  inv U319 ( .a(n318), .out(\sig_prgm_register/or_signal [317]) );
  inv U320 ( .a(n319), .out(\sig_prgm_register/or_signal [318]) );
  inv U321 ( .a(n320), .out(\sig_prgm_register/or_signal [319]) );
  inv U322 ( .a(n321), .out(\sig_prgm_register/or_signal [320]) );
  inv U323 ( .a(n322), .out(\sig_prgm_register/or_signal [321]) );
  inv U324 ( .a(n323), .out(\sig_prgm_register/or_signal [322]) );
  inv U325 ( .a(n324), .out(\sig_prgm_register/or_signal [323]) );
  inv U326 ( .a(n325), .out(\sig_prgm_register/or_signal [324]) );
  inv U327 ( .a(n326), .out(\sig_prgm_register/or_signal [325]) );
  inv U328 ( .a(n327), .out(\sig_prgm_register/or_signal [326]) );
  inv U329 ( .a(n328), .out(\sig_prgm_register/or_signal [327]) );
  inv U330 ( .a(n329), .out(\sig_prgm_register/or_signal [328]) );
  inv U331 ( .a(n330), .out(\sig_prgm_register/or_signal [329]) );
  inv U332 ( .a(n331), .out(\sig_prgm_register/or_signal [330]) );
  inv U333 ( .a(n332), .out(\sig_prgm_register/or_signal [331]) );
  inv U334 ( .a(n333), .out(\sig_prgm_register/or_signal [332]) );
  inv U335 ( .a(n334), .out(\sig_prgm_register/or_signal [333]) );
  inv U336 ( .a(n335), .out(\sig_prgm_register/or_signal [334]) );
  inv U337 ( .a(n336), .out(\sig_prgm_register/or_signal [335]) );
  inv U338 ( .a(n337), .out(\sig_prgm_register/or_signal [336]) );
  inv U339 ( .a(n338), .out(\sig_prgm_register/or_signal [337]) );
  inv U340 ( .a(n339), .out(\sig_prgm_register/or_signal [338]) );
  inv U341 ( .a(n340), .out(\sig_prgm_register/or_signal [339]) );
  inv U342 ( .a(n341), .out(\sig_prgm_register/or_signal [340]) );
  inv U343 ( .a(n342), .out(\sig_prgm_register/or_signal [341]) );
  inv U344 ( .a(n343), .out(\sig_prgm_register/or_signal [342]) );
  inv U345 ( .a(n344), .out(\sig_prgm_register/or_signal [343]) );
  inv U346 ( .a(n345), .out(\sig_prgm_register/or_signal [344]) );
  inv U347 ( .a(n346), .out(\sig_prgm_register/or_signal [345]) );
  inv U348 ( .a(n347), .out(\sig_prgm_register/or_signal [346]) );
  inv U349 ( .a(n348), .out(\sig_prgm_register/or_signal [347]) );
  inv U350 ( .a(n349), .out(\sig_prgm_register/or_signal [348]) );
  inv U351 ( .a(n350), .out(\sig_prgm_register/or_signal [349]) );
  inv U352 ( .a(n351), .out(\sig_prgm_register/or_signal [350]) );
  inv U353 ( .a(n352), .out(\sig_prgm_register/or_signal [351]) );
  inv U354 ( .a(n353), .out(\sig_prgm_register/or_signal [352]) );
  inv U355 ( .a(n354), .out(\sig_prgm_register/or_signal [353]) );
  inv U356 ( .a(n355), .out(\sig_prgm_register/or_signal [354]) );
  inv U357 ( .a(n356), .out(\sig_prgm_register/or_signal [355]) );
  inv U358 ( .a(n357), .out(\sig_prgm_register/or_signal [356]) );
  inv U359 ( .a(n358), .out(\sig_prgm_register/or_signal [357]) );
  inv U360 ( .a(n359), .out(\sig_prgm_register/or_signal [358]) );
  inv U361 ( .a(n360), .out(\sig_prgm_register/or_signal [359]) );
  inv U362 ( .a(n361), .out(\sig_prgm_register/or_signal [360]) );
  inv U363 ( .a(n362), .out(\sig_prgm_register/or_signal [361]) );
  inv U364 ( .a(n363), .out(\sig_prgm_register/or_signal [362]) );
  inv U365 ( .a(n364), .out(\sig_prgm_register/or_signal [363]) );
  inv U366 ( .a(n365), .out(\sig_prgm_register/or_signal [364]) );
  inv U367 ( .a(n366), .out(\sig_prgm_register/or_signal [365]) );
  inv U368 ( .a(n367), .out(\sig_prgm_register/or_signal [366]) );
  inv U369 ( .a(n368), .out(\sig_prgm_register/or_signal [367]) );
  inv U370 ( .a(n369), .out(\sig_prgm_register/or_signal [368]) );
  inv U371 ( .a(n370), .out(\sig_prgm_register/or_signal [369]) );
  inv U372 ( .a(n371), .out(\sig_prgm_register/or_signal [370]) );
  inv U373 ( .a(n372), .out(\sig_prgm_register/or_signal [371]) );
  inv U374 ( .a(n373), .out(\sig_prgm_register/or_signal [372]) );
  inv U375 ( .a(n374), .out(\sig_prgm_register/or_signal [373]) );
  inv U376 ( .a(n375), .out(\sig_prgm_register/or_signal [374]) );
  inv U377 ( .a(n376), .out(\sig_prgm_register/or_signal [375]) );
  inv U378 ( .a(n377), .out(\sig_prgm_register/or_signal [376]) );
  inv U379 ( .a(n378), .out(\sig_prgm_register/or_signal [377]) );
  inv U380 ( .a(n379), .out(\sig_prgm_register/or_signal [378]) );
  inv U381 ( .a(n380), .out(\sig_prgm_register/or_signal [379]) );
  inv U382 ( .a(n381), .out(\sig_prgm_register/or_signal [380]) );
  inv U383 ( .a(n382), .out(\sig_prgm_register/or_signal [381]) );
  inv U384 ( .a(n383), .out(\sig_prgm_register/or_signal [382]) );
  inv U385 ( .a(n384), .out(\sig_prgm_register/or_signal [383]) );
  inv U386 ( .a(n385), .out(\sig_prgm_register/or_signal [384]) );
  inv U387 ( .a(n386), .out(\sig_prgm_register/or_signal [385]) );
  inv U388 ( .a(n387), .out(\sig_prgm_register/or_signal [386]) );
  inv U389 ( .a(n388), .out(\sig_prgm_register/or_signal [387]) );
  inv U390 ( .a(n389), .out(\sig_prgm_register/or_signal [388]) );
  inv U391 ( .a(n390), .out(\sig_prgm_register/or_signal [389]) );
  inv U392 ( .a(n391), .out(\sig_prgm_register/or_signal [390]) );
  inv U393 ( .a(n392), .out(\sig_prgm_register/or_signal [391]) );
  inv U394 ( .a(n393), .out(\sig_prgm_register/or_signal [392]) );
  inv U395 ( .a(n394), .out(\sig_prgm_register/or_signal [393]) );
  inv U396 ( .a(n395), .out(\sig_prgm_register/or_signal [394]) );
  inv U397 ( .a(n396), .out(\sig_prgm_register/or_signal [395]) );
  inv U398 ( .a(n397), .out(\sig_prgm_register/or_signal [396]) );
  inv U399 ( .a(n398), .out(\sig_prgm_register/or_signal [397]) );
  inv U400 ( .a(n399), .out(\sig_prgm_register/or_signal [398]) );
  inv U401 ( .a(n400), .out(\sig_prgm_register/or_signal [399]) );
  inv U402 ( .a(n401), .out(\sig_prgm_register/or_signal [400]) );
  inv U403 ( .a(n402), .out(\sig_prgm_register/or_signal [401]) );
  inv U404 ( .a(n403), .out(\sig_prgm_register/or_signal [402]) );
  inv U405 ( .a(n404), .out(\sig_prgm_register/or_signal [403]) );
  inv U406 ( .a(n405), .out(\sig_prgm_register/or_signal [404]) );
  inv U407 ( .a(n406), .out(\sig_prgm_register/or_signal [405]) );
  inv U408 ( .a(n407), .out(\sig_prgm_register/or_signal [406]) );
  inv U409 ( .a(n408), .out(\sig_prgm_register/or_signal [407]) );
  inv U410 ( .a(n409), .out(\sig_prgm_register/or_signal [408]) );
  inv U411 ( .a(n410), .out(\sig_prgm_register/or_signal [409]) );
  inv U412 ( .a(n411), .out(\sig_prgm_register/or_signal [410]) );
  inv U413 ( .a(n412), .out(\sig_prgm_register/or_signal [411]) );
  inv U414 ( .a(n413), .out(\sig_prgm_register/or_signal [412]) );
  inv U415 ( .a(n414), .out(\sig_prgm_register/or_signal [413]) );
  inv U416 ( .a(n415), .out(\sig_prgm_register/or_signal [414]) );
  inv U417 ( .a(n416), .out(\sig_prgm_register/or_signal [415]) );
  inv U418 ( .a(n417), .out(\sig_prgm_register/or_signal [416]) );
  inv U419 ( .a(n418), .out(\sig_prgm_register/or_signal [417]) );
  inv U420 ( .a(n419), .out(\sig_prgm_register/or_signal [418]) );
  inv U421 ( .a(n420), .out(\sig_prgm_register/or_signal [419]) );
  inv U422 ( .a(n421), .out(\sig_prgm_register/or_signal [420]) );
  inv U423 ( .a(n422), .out(\sig_prgm_register/or_signal [421]) );
  inv U424 ( .a(n423), .out(\sig_prgm_register/or_signal [422]) );
  inv U425 ( .a(n424), .out(\sig_prgm_register/or_signal [423]) );
  inv U426 ( .a(n425), .out(\sig_prgm_register/or_signal [424]) );
  inv U427 ( .a(n426), .out(\sig_prgm_register/or_signal [425]) );
  inv U428 ( .a(n427), .out(\sig_prgm_register/or_signal [426]) );
  inv U429 ( .a(n428), .out(\sig_prgm_register/or_signal [427]) );
  inv U430 ( .a(n429), .out(\sig_prgm_register/or_signal [428]) );
  inv U431 ( .a(n430), .out(\sig_prgm_register/or_signal [429]) );
  inv U432 ( .a(n431), .out(\sig_prgm_register/or_signal [430]) );
  inv U433 ( .a(n432), .out(\sig_prgm_register/or_signal [431]) );
  inv U434 ( .a(n433), .out(\sig_prgm_register/or_signal [432]) );
  inv U435 ( .a(n434), .out(\sig_prgm_register/or_signal [433]) );
  inv U436 ( .a(n435), .out(\sig_prgm_register/or_signal [434]) );
  inv U437 ( .a(n436), .out(\sig_prgm_register/or_signal [435]) );
  inv U438 ( .a(n437), .out(\sig_prgm_register/or_signal [436]) );
  inv U439 ( .a(n438), .out(\sig_prgm_register/or_signal [437]) );
  inv U440 ( .a(n439), .out(\sig_prgm_register/or_signal [438]) );
  inv U441 ( .a(n440), .out(\sig_prgm_register/or_signal [439]) );
  inv U442 ( .a(n441), .out(\sig_prgm_register/or_signal [440]) );
  inv U443 ( .a(n442), .out(\sig_prgm_register/or_signal [441]) );
  inv U444 ( .a(n443), .out(\sig_prgm_register/or_signal [442]) );
  inv U445 ( .a(n444), .out(\sig_prgm_register/or_signal [443]) );
  inv U446 ( .a(n445), .out(\sig_prgm_register/or_signal [444]) );
  inv U447 ( .a(n446), .out(\sig_prgm_register/or_signal [445]) );
  inv U448 ( .a(n447), .out(\sig_prgm_register/or_signal [446]) );
  inv U449 ( .a(n448), .out(\sig_prgm_register/or_signal [447]) );
  inv U450 ( .a(n449), .out(\sig_prgm_register/or_signal [448]) );
  inv U451 ( .a(n450), .out(\sig_prgm_register/or_signal [449]) );
  inv U452 ( .a(n451), .out(\sig_prgm_register/or_signal [450]) );
  inv U453 ( .a(n452), .out(\sig_prgm_register/or_signal [451]) );
  inv U454 ( .a(n453), .out(\sig_prgm_register/or_signal [452]) );
  inv U455 ( .a(n454), .out(\sig_prgm_register/or_signal [453]) );
  inv U456 ( .a(n455), .out(\sig_prgm_register/or_signal [454]) );
  inv U457 ( .a(n456), .out(\sig_prgm_register/or_signal [455]) );
  inv U458 ( .a(n457), .out(\sig_prgm_register/or_signal [456]) );
  inv U459 ( .a(n458), .out(\sig_prgm_register/or_signal [457]) );
  inv U460 ( .a(n459), .out(\sig_prgm_register/or_signal [458]) );
  inv U461 ( .a(n460), .out(\sig_prgm_register/or_signal [459]) );
  inv U462 ( .a(n461), .out(\sig_prgm_register/or_signal [460]) );
  inv U463 ( .a(n462), .out(\sig_prgm_register/or_signal [461]) );
  inv U464 ( .a(n463), .out(\sig_prgm_register/or_signal [462]) );
  inv U465 ( .a(n464), .out(\sig_prgm_register/or_signal [463]) );
  inv U466 ( .a(n465), .out(\sig_prgm_register/or_signal [464]) );
  inv U467 ( .a(n466), .out(\sig_prgm_register/or_signal [465]) );
  inv U468 ( .a(n467), .out(\sig_prgm_register/or_signal [466]) );
  inv U469 ( .a(n468), .out(\sig_prgm_register/or_signal [467]) );
  inv U470 ( .a(n469), .out(\sig_prgm_register/or_signal [468]) );
  inv U471 ( .a(n470), .out(\sig_prgm_register/or_signal [469]) );
  inv U472 ( .a(n471), .out(\sig_prgm_register/or_signal [470]) );
  inv U473 ( .a(n472), .out(\sig_prgm_register/or_signal [471]) );
  inv U474 ( .a(n473), .out(\sig_prgm_register/or_signal [472]) );
  inv U475 ( .a(n474), .out(\sig_prgm_register/or_signal [473]) );
  inv U476 ( .a(n475), .out(\sig_prgm_register/or_signal [474]) );
  inv U477 ( .a(n476), .out(\sig_prgm_register/or_signal [475]) );
  inv U478 ( .a(n477), .out(\sig_prgm_register/or_signal [476]) );
  inv U479 ( .a(n478), .out(\sig_prgm_register/or_signal [477]) );
  inv U480 ( .a(n479), .out(\sig_prgm_register/or_signal [478]) );
  inv U481 ( .a(n480), .out(\sig_prgm_register/or_signal [479]) );
  inv U482 ( .a(n481), .out(\sig_prgm_register/or_signal [480]) );
  inv U483 ( .a(n482), .out(\sig_prgm_register/or_signal [481]) );
  inv U484 ( .a(n483), .out(\sig_prgm_register/or_signal [482]) );
  inv U485 ( .a(n484), .out(\sig_prgm_register/or_signal [483]) );
  inv U486 ( .a(n485), .out(\sig_prgm_register/or_signal [484]) );
  inv U487 ( .a(n486), .out(\sig_prgm_register/or_signal [485]) );
  inv U488 ( .a(n487), .out(\sig_prgm_register/or_signal [486]) );
  inv U489 ( .a(n488), .out(\sig_prgm_register/or_signal [487]) );
  inv U490 ( .a(n489), .out(\sig_prgm_register/or_signal [488]) );
  inv U491 ( .a(n490), .out(\sig_prgm_register/or_signal [489]) );
  inv U492 ( .a(n491), .out(\sig_prgm_register/or_signal [490]) );
  inv U493 ( .a(n492), .out(\sig_prgm_register/or_signal [491]) );
  inv U494 ( .a(n493), .out(\sig_prgm_register/or_signal [492]) );
  inv U495 ( .a(n494), .out(\sig_prgm_register/or_signal [493]) );
  inv U496 ( .a(n495), .out(\sig_prgm_register/or_signal [494]) );
  inv U497 ( .a(n496), .out(\sig_prgm_register/or_signal [495]) );
  inv U498 ( .a(n497), .out(\sig_prgm_register/or_signal [496]) );
  inv U499 ( .a(n498), .out(\sig_prgm_register/or_signal [497]) );
  inv U500 ( .a(n499), .out(\sig_prgm_register/or_signal [498]) );
  inv U501 ( .a(n500), .out(\sig_prgm_register/or_signal [499]) );
  inv U502 ( .a(n501), .out(\sig_prgm_register/or_signal [500]) );
  inv U503 ( .a(n502), .out(\sig_prgm_register/or_signal [501]) );
  inv U504 ( .a(n503), .out(\sig_prgm_register/or_signal [502]) );
  inv U505 ( .a(n504), .out(\sig_prgm_register/or_signal [503]) );
  inv U506 ( .a(n505), .out(\sig_prgm_register/or_signal [504]) );
  inv U507 ( .a(n506), .out(\sig_prgm_register/or_signal [505]) );
  inv U508 ( .a(n507), .out(\sig_prgm_register/or_signal [506]) );
  inv U509 ( .a(n508), .out(\sig_prgm_register/or_signal [507]) );
  inv U510 ( .a(n509), .out(\sig_prgm_register/or_signal [508]) );
  inv U511 ( .a(n510), .out(\sig_prgm_register/or_signal [509]) );
  inv U512 ( .a(n511), .out(\sig_prgm_register/or_signal [510]) );
  inv U513 ( .a(n512), .out(\sig_prgm_register/or_signal [511]) );
  inv U514 ( .a(n513), .out(\sig_prgm_register/or_signal [512]) );
  inv U515 ( .a(n514), .out(\sig_prgm_register/or_signal [513]) );
  inv U516 ( .a(n515), .out(\sig_prgm_register/or_signal [514]) );
  inv U517 ( .a(n516), .out(\sig_prgm_register/or_signal [515]) );
  inv U518 ( .a(n517), .out(\sig_prgm_register/or_signal [516]) );
  inv U519 ( .a(n518), .out(\sig_prgm_register/or_signal [517]) );
  inv U520 ( .a(n519), .out(\sig_prgm_register/or_signal [518]) );
  inv U521 ( .a(n520), .out(\sig_prgm_register/or_signal [519]) );
  inv U522 ( .a(n521), .out(\sig_prgm_register/or_signal [520]) );
  inv U523 ( .a(n522), .out(\sig_prgm_register/or_signal [521]) );
  inv U524 ( .a(n523), .out(\sig_prgm_register/or_signal [522]) );
  inv U525 ( .a(n524), .out(\sig_prgm_register/or_signal [523]) );
  inv U526 ( .a(n525), .out(\sig_prgm_register/or_signal [524]) );
  inv U527 ( .a(n526), .out(\sig_prgm_register/or_signal [525]) );
  inv U528 ( .a(n527), .out(\sig_prgm_register/or_signal [526]) );
  inv U529 ( .a(n528), .out(\sig_prgm_register/or_signal [527]) );
  inv U530 ( .a(n529), .out(\sig_prgm_register/or_signal [528]) );
  inv U531 ( .a(n530), .out(\sig_prgm_register/or_signal [529]) );
  inv U532 ( .a(n531), .out(\sig_prgm_register/or_signal [530]) );
  inv U533 ( .a(n532), .out(\sig_prgm_register/or_signal [531]) );
  inv U534 ( .a(n533), .out(\sig_prgm_register/or_signal [532]) );
  inv U535 ( .a(n534), .out(\sig_prgm_register/or_signal [533]) );
  inv U536 ( .a(n535), .out(\sig_prgm_register/or_signal [534]) );
  inv U537 ( .a(n536), .out(\sig_prgm_register/or_signal [535]) );
  inv U538 ( .a(n537), .out(\sig_prgm_register/or_signal [536]) );
  inv U539 ( .a(n538), .out(\sig_prgm_register/or_signal [537]) );
  inv U540 ( .a(n539), .out(\sig_prgm_register/or_signal [538]) );
  inv U541 ( .a(n540), .out(\sig_prgm_register/or_signal [539]) );
  inv U542 ( .a(n541), .out(\sig_prgm_register/or_signal [540]) );
  inv U543 ( .a(n542), .out(\sig_prgm_register/or_signal [541]) );
  inv U544 ( .a(n543), .out(\sig_prgm_register/or_signal [542]) );
  inv U545 ( .a(n544), .out(\sig_prgm_register/or_signal [543]) );
  inv U546 ( .a(n545), .out(\sig_prgm_register/or_signal [544]) );
  inv U547 ( .a(n546), .out(\sig_prgm_register/or_signal [545]) );
  inv U548 ( .a(n547), .out(\sig_prgm_register/or_signal [546]) );
  inv U549 ( .a(n548), .out(\sig_prgm_register/or_signal [547]) );
  inv U550 ( .a(n549), .out(\sig_prgm_register/or_signal [548]) );
  inv U551 ( .a(n550), .out(\sig_prgm_register/or_signal [549]) );
  inv U552 ( .a(n551), .out(\sig_prgm_register/or_signal [550]) );
  inv U553 ( .a(n552), .out(\sig_prgm_register/or_signal [551]) );
  inv U554 ( .a(n553), .out(\sig_prgm_register/or_signal [552]) );
  inv U555 ( .a(n554), .out(\sig_prgm_register/or_signal [553]) );
  inv U556 ( .a(n555), .out(\sig_prgm_register/or_signal [554]) );
  inv U557 ( .a(n556), .out(\sig_prgm_register/or_signal [555]) );
  inv U558 ( .a(n557), .out(\sig_prgm_register/or_signal [556]) );
  inv U559 ( .a(n558), .out(\sig_prgm_register/or_signal [557]) );
  inv U560 ( .a(n559), .out(\sig_prgm_register/or_signal [558]) );
  inv U561 ( .a(n560), .out(\sig_prgm_register/or_signal [559]) );
  inv U562 ( .a(n561), .out(\sig_prgm_register/or_signal [560]) );
  inv U563 ( .a(n562), .out(\sig_prgm_register/or_signal [561]) );
  inv U564 ( .a(n563), .out(\sig_prgm_register/or_signal [562]) );
  inv U565 ( .a(n564), .out(\sig_prgm_register/or_signal [563]) );
  inv U566 ( .a(n565), .out(\sig_prgm_register/or_signal [564]) );
  inv U567 ( .a(n566), .out(\sig_prgm_register/or_signal [565]) );
  inv U568 ( .a(n567), .out(\sig_prgm_register/or_signal [566]) );
  inv U569 ( .a(n568), .out(\sig_prgm_register/or_signal [567]) );
  inv U570 ( .a(n569), .out(\sig_prgm_register/or_signal [568]) );
  inv U571 ( .a(n570), .out(\sig_prgm_register/or_signal [569]) );
  inv U572 ( .a(n571), .out(\sig_prgm_register/or_signal [570]) );
  inv U573 ( .a(n572), .out(\sig_prgm_register/or_signal [571]) );
  inv U574 ( .a(n573), .out(\sig_prgm_register/or_signal [572]) );
  inv U575 ( .a(n574), .out(\sig_prgm_register/or_signal [573]) );
  inv U576 ( .a(n575), .out(\sig_prgm_register/or_signal [574]) );
  inv U577 ( .a(n576), .out(\sig_prgm_register/or_signal [575]) );
  inv U578 ( .a(n577), .out(\sig_prgm_register/or_signal [576]) );
  inv U579 ( .a(n578), .out(\sig_prgm_register/or_signal [577]) );
  inv U580 ( .a(n579), .out(\sig_prgm_register/or_signal [578]) );
  inv U581 ( .a(n580), .out(\sig_prgm_register/or_signal [579]) );
  inv U582 ( .a(n581), .out(\sig_prgm_register/or_signal [580]) );
  inv U583 ( .a(n582), .out(\sig_prgm_register/or_signal [581]) );
  inv U584 ( .a(n583), .out(\sig_prgm_register/or_signal [582]) );
  inv U585 ( .a(n584), .out(\sig_prgm_register/or_signal [583]) );
  inv U586 ( .a(n585), .out(\sig_prgm_register/or_signal [584]) );
  inv U587 ( .a(n586), .out(\sig_prgm_register/or_signal [585]) );
  inv U588 ( .a(n587), .out(\sig_prgm_register/or_signal [586]) );
  inv U589 ( .a(n588), .out(\sig_prgm_register/or_signal [587]) );
  inv U590 ( .a(n589), .out(\sig_prgm_register/or_signal [588]) );
  inv U591 ( .a(n590), .out(\sig_prgm_register/or_signal [589]) );
  inv U592 ( .a(n591), .out(\sig_prgm_register/or_signal [590]) );
  inv U593 ( .a(n592), .out(\sig_prgm_register/or_signal [591]) );
  inv U594 ( .a(n593), .out(\sig_prgm_register/or_signal [592]) );
  inv U595 ( .a(n594), .out(\sig_prgm_register/or_signal [593]) );
  inv U596 ( .a(n595), .out(\sig_prgm_register/or_signal [594]) );
  inv U597 ( .a(n596), .out(\sig_prgm_register/or_signal [595]) );
  inv U598 ( .a(n597), .out(\sig_prgm_register/or_signal [596]) );
  inv U599 ( .a(n598), .out(\sig_prgm_register/or_signal [597]) );
  inv U600 ( .a(n599), .out(\sig_prgm_register/or_signal [598]) );
  inv U601 ( .a(n600), .out(\sig_prgm_register/or_signal [599]) );
  inv U602 ( .a(n601), .out(\sig_prgm_register/or_signal [600]) );
  inv U603 ( .a(n602), .out(\sig_prgm_register/or_signal [601]) );
  inv U604 ( .a(n603), .out(\sig_prgm_register/or_signal [602]) );
  inv U605 ( .a(n604), .out(\sig_prgm_register/or_signal [603]) );
  inv U606 ( .a(n605), .out(\sig_prgm_register/or_signal [604]) );
  inv U607 ( .a(n606), .out(\sig_prgm_register/or_signal [605]) );
  inv U608 ( .a(n607), .out(\sig_prgm_register/or_signal [606]) );
  inv U609 ( .a(n608), .out(\sig_prgm_register/or_signal [607]) );
  inv U610 ( .a(n609), .out(\sig_prgm_register/or_signal [608]) );
  inv U611 ( .a(n610), .out(\sig_prgm_register/or_signal [609]) );
  inv U612 ( .a(n611), .out(\sig_prgm_register/or_signal [610]) );
  inv U613 ( .a(n612), .out(\sig_prgm_register/or_signal [611]) );
  inv U614 ( .a(n613), .out(\sig_prgm_register/or_signal [612]) );
  inv U615 ( .a(n614), .out(\sig_prgm_register/or_signal [613]) );
  inv U616 ( .a(n615), .out(\sig_prgm_register/or_signal [614]) );
  inv U617 ( .a(n616), .out(\sig_prgm_register/or_signal [615]) );
  inv U618 ( .a(n617), .out(\sig_prgm_register/or_signal [616]) );
  inv U619 ( .a(n618), .out(\sig_prgm_register/or_signal [617]) );
  inv U620 ( .a(n619), .out(\sig_prgm_register/or_signal [618]) );
  inv U621 ( .a(n620), .out(\sig_prgm_register/or_signal [619]) );
  inv U622 ( .a(n621), .out(\sig_prgm_register/or_signal [620]) );
  inv U623 ( .a(n622), .out(\sig_prgm_register/or_signal [621]) );
  inv U624 ( .a(n623), .out(\sig_prgm_register/or_signal [622]) );
  inv U625 ( .a(n624), .out(\sig_prgm_register/or_signal [623]) );
  inv U626 ( .a(n625), .out(\sig_prgm_register/or_signal [624]) );
  inv U627 ( .a(n626), .out(\sig_prgm_register/or_signal [625]) );
  inv U628 ( .a(n627), .out(\sig_prgm_register/or_signal [626]) );
  inv U629 ( .a(n628), .out(\sig_prgm_register/or_signal [627]) );
  inv U630 ( .a(n629), .out(\sig_prgm_register/or_signal [628]) );
  inv U631 ( .a(n630), .out(\sig_prgm_register/or_signal [629]) );
  inv U632 ( .a(n631), .out(\sig_prgm_register/or_signal [630]) );
  inv U633 ( .a(n632), .out(\sig_prgm_register/or_signal [631]) );
  inv U634 ( .a(n633), .out(\sig_prgm_register/or_signal [632]) );
  inv U635 ( .a(n634), .out(\sig_prgm_register/or_signal [633]) );
  inv U636 ( .a(n635), .out(\sig_prgm_register/or_signal [634]) );
  inv U637 ( .a(n636), .out(\sig_prgm_register/or_signal [635]) );
  inv U638 ( .a(n637), .out(\sig_prgm_register/or_signal [636]) );
  inv U639 ( .a(n638), .out(\sig_prgm_register/or_signal [637]) );
  inv U640 ( .a(n639), .out(\sig_prgm_register/or_signal [638]) );
  inv U641 ( .a(n640), .out(\sig_prgm_register/or_signal [639]) );
  inv U642 ( .a(n641), .out(\sig_prgm_register/or_signal [640]) );
  inv U643 ( .a(n642), .out(\sig_prgm_register/or_signal [641]) );
  inv U644 ( .a(n643), .out(\sig_prgm_register/or_signal [642]) );
  inv U645 ( .a(n644), .out(\sig_prgm_register/or_signal [643]) );
  inv U646 ( .a(n645), .out(\sig_prgm_register/or_signal [644]) );
  inv U647 ( .a(n646), .out(\sig_prgm_register/or_signal [645]) );
  inv U648 ( .a(n647), .out(\sig_prgm_register/or_signal [646]) );
  inv U649 ( .a(n648), .out(\sig_prgm_register/or_signal [647]) );
  inv U650 ( .a(n649), .out(\sig_prgm_register/or_signal [648]) );
  inv U651 ( .a(n650), .out(\sig_prgm_register/or_signal [649]) );
  inv U652 ( .a(n651), .out(\sig_prgm_register/or_signal [650]) );
  inv U653 ( .a(n652), .out(\sig_prgm_register/or_signal [651]) );
  inv U654 ( .a(n653), .out(\sig_prgm_register/or_signal [652]) );
  inv U655 ( .a(n654), .out(\sig_prgm_register/or_signal [653]) );
  inv U656 ( .a(n655), .out(\sig_prgm_register/or_signal [654]) );
  inv U657 ( .a(n656), .out(\sig_prgm_register/or_signal [655]) );
  inv U658 ( .a(n657), .out(\sig_prgm_register/or_signal [656]) );
  inv U659 ( .a(n658), .out(\sig_prgm_register/or_signal [657]) );
  inv U660 ( .a(n659), .out(\sig_prgm_register/or_signal [658]) );
  inv U661 ( .a(n660), .out(\sig_prgm_register/or_signal [659]) );
  inv U662 ( .a(n661), .out(\sig_prgm_register/or_signal [660]) );
  inv U663 ( .a(n662), .out(\sig_prgm_register/or_signal [661]) );
  inv U664 ( .a(n663), .out(\sig_prgm_register/or_signal [662]) );
  inv U665 ( .a(n664), .out(\sig_prgm_register/or_signal [663]) );
  inv U666 ( .a(n665), .out(\sig_prgm_register/or_signal [664]) );
  inv U667 ( .a(n666), .out(\sig_prgm_register/or_signal [665]) );
  inv U668 ( .a(n667), .out(\sig_prgm_register/or_signal [666]) );
  inv U669 ( .a(n668), .out(\sig_prgm_register/or_signal [667]) );
  inv U670 ( .a(n669), .out(\sig_prgm_register/or_signal [668]) );
  inv U671 ( .a(n670), .out(\sig_prgm_register/or_signal [669]) );
  inv U672 ( .a(n671), .out(\sig_prgm_register/or_signal [670]) );
  inv U673 ( .a(n672), .out(\sig_prgm_register/or_signal [671]) );
  inv U674 ( .a(n673), .out(\sig_prgm_register/or_signal [672]) );
  inv U675 ( .a(n674), .out(\sig_prgm_register/or_signal [673]) );
  inv U676 ( .a(n675), .out(\sig_prgm_register/or_signal [674]) );
  inv U677 ( .a(n676), .out(\sig_prgm_register/or_signal [675]) );
  inv U678 ( .a(n677), .out(\sig_prgm_register/or_signal [676]) );
  inv U679 ( .a(n678), .out(\sig_prgm_register/or_signal [677]) );
  inv U680 ( .a(n679), .out(\sig_prgm_register/or_signal [678]) );
  inv U681 ( .a(n680), .out(\sig_prgm_register/or_signal [679]) );
  inv U682 ( .a(n681), .out(\sig_prgm_register/or_signal [680]) );
  inv U683 ( .a(n682), .out(\sig_prgm_register/or_signal [681]) );
  inv U684 ( .a(n683), .out(\sig_prgm_register/or_signal [682]) );
  inv U685 ( .a(n684), .out(\sig_prgm_register/or_signal [683]) );
  inv U686 ( .a(n685), .out(\sig_prgm_register/or_signal [684]) );
  inv U687 ( .a(n686), .out(\sig_prgm_register/or_signal [685]) );
  inv U688 ( .a(n687), .out(\sig_prgm_register/or_signal [686]) );
  inv U689 ( .a(n688), .out(\sig_prgm_register/or_signal [687]) );
  inv U690 ( .a(n689), .out(\sig_prgm_register/or_signal [688]) );
  inv U691 ( .a(n690), .out(\sig_prgm_register/or_signal [689]) );
  inv U692 ( .a(n691), .out(\sig_prgm_register/or_signal [690]) );
  inv U693 ( .a(n692), .out(\sig_prgm_register/or_signal [691]) );
  inv U694 ( .a(n693), .out(\sig_prgm_register/or_signal [692]) );
  inv U695 ( .a(n694), .out(\sig_prgm_register/or_signal [693]) );
  inv U696 ( .a(n695), .out(\sig_prgm_register/or_signal [694]) );
  inv U697 ( .a(n696), .out(\sig_prgm_register/or_signal [695]) );
  inv U698 ( .a(n697), .out(\sig_prgm_register/or_signal [696]) );
  inv U699 ( .a(n698), .out(\sig_prgm_register/or_signal [697]) );
  inv U700 ( .a(n699), .out(\sig_prgm_register/or_signal [698]) );
  inv U701 ( .a(n700), .out(\sig_prgm_register/or_signal [699]) );
  inv U702 ( .a(n701), .out(\sig_prgm_register/or_signal [700]) );
  inv U703 ( .a(n702), .out(\sig_prgm_register/or_signal [701]) );
  inv U704 ( .a(n703), .out(\sig_prgm_register/or_signal [702]) );
  inv U705 ( .a(n704), .out(\sig_prgm_register/or_signal [703]) );
  inv U706 ( .a(n705), .out(\sig_prgm_register/or_signal [704]) );
  inv U707 ( .a(n706), .out(\sig_prgm_register/or_signal [705]) );
  inv U708 ( .a(n707), .out(\sig_prgm_register/or_signal [706]) );
  inv U709 ( .a(n708), .out(\sig_prgm_register/or_signal [707]) );
  inv U710 ( .a(n709), .out(\sig_prgm_register/or_signal [708]) );
  inv U711 ( .a(n710), .out(\sig_prgm_register/or_signal [709]) );
  inv U712 ( .a(n711), .out(\sig_prgm_register/or_signal [710]) );
  inv U713 ( .a(n712), .out(\sig_prgm_register/or_signal [711]) );
  inv U714 ( .a(n713), .out(\sig_prgm_register/or_signal [712]) );
  inv U715 ( .a(n714), .out(\sig_prgm_register/or_signal [713]) );
  inv U716 ( .a(n715), .out(\sig_prgm_register/or_signal [714]) );
  inv U717 ( .a(n716), .out(\sig_prgm_register/or_signal [715]) );
  inv U718 ( .a(n717), .out(\sig_prgm_register/or_signal [716]) );
  inv U719 ( .a(n718), .out(\sig_prgm_register/or_signal [717]) );
  inv U720 ( .a(n719), .out(\sig_prgm_register/or_signal [718]) );
  inv U721 ( .a(n720), .out(\sig_prgm_register/or_signal [719]) );
  inv U722 ( .a(n721), .out(\sig_prgm_register/or_signal [720]) );
  inv U723 ( .a(n722), .out(\sig_prgm_register/or_signal [721]) );
  inv U724 ( .a(n723), .out(\sig_prgm_register/or_signal [722]) );
  inv U725 ( .a(n724), .out(\sig_prgm_register/or_signal [723]) );
  inv U726 ( .a(n725), .out(\sig_prgm_register/or_signal [724]) );
  inv U727 ( .a(n726), .out(\sig_prgm_register/or_signal [725]) );
  inv U728 ( .a(n727), .out(\sig_prgm_register/or_signal [726]) );
  inv U729 ( .a(n728), .out(\sig_prgm_register/or_signal [727]) );
  inv U730 ( .a(n729), .out(\sig_prgm_register/or_signal [728]) );
  inv U731 ( .a(n730), .out(\sig_prgm_register/or_signal [729]) );
  inv U732 ( .a(n731), .out(\sig_prgm_register/or_signal [730]) );
  inv U733 ( .a(n732), .out(\sig_prgm_register/or_signal [731]) );
  inv U734 ( .a(n733), .out(\sig_prgm_register/or_signal [732]) );
  inv U735 ( .a(n734), .out(\sig_prgm_register/or_signal [733]) );
  inv U736 ( .a(n735), .out(\sig_prgm_register/or_signal [734]) );
  inv U737 ( .a(n736), .out(\sig_prgm_register/or_signal [735]) );
  inv U738 ( .a(n737), .out(\sig_prgm_register/or_signal [736]) );
  inv U739 ( .a(n738), .out(\sig_prgm_register/or_signal [737]) );
  inv U740 ( .a(n739), .out(\sig_prgm_register/or_signal [738]) );
  inv U741 ( .a(n740), .out(\sig_prgm_register/or_signal [739]) );
  inv U742 ( .a(n741), .out(\sig_prgm_register/or_signal [740]) );
  inv U743 ( .a(n742), .out(\sig_prgm_register/or_signal [741]) );
  inv U744 ( .a(n743), .out(\sig_prgm_register/or_signal [742]) );
  inv U745 ( .a(n744), .out(\sig_prgm_register/or_signal [743]) );
  inv U746 ( .a(n745), .out(\sig_prgm_register/or_signal [744]) );
  inv U747 ( .a(n746), .out(\sig_prgm_register/or_signal [745]) );
  inv U748 ( .a(n747), .out(\sig_prgm_register/or_signal [746]) );
  inv U749 ( .a(n748), .out(\sig_prgm_register/or_signal [747]) );
  inv U750 ( .a(n749), .out(\sig_prgm_register/or_signal [748]) );
  inv U751 ( .a(n750), .out(\sig_prgm_register/or_signal [749]) );
  inv U752 ( .a(n751), .out(\sig_prgm_register/or_signal [750]) );
  inv U753 ( .a(n752), .out(\sig_prgm_register/or_signal [751]) );
  inv U754 ( .a(n753), .out(\sig_prgm_register/or_signal [752]) );
  inv U755 ( .a(n754), .out(\sig_prgm_register/or_signal [753]) );
  inv U756 ( .a(n755), .out(\sig_prgm_register/or_signal [754]) );
  inv U757 ( .a(n756), .out(\sig_prgm_register/or_signal [755]) );
  inv U758 ( .a(n757), .out(\sig_prgm_register/or_signal [756]) );
  inv U759 ( .a(n758), .out(\sig_prgm_register/or_signal [757]) );
  inv U760 ( .a(n759), .out(\sig_prgm_register/or_signal [758]) );
  inv U761 ( .a(n760), .out(\sig_prgm_register/or_signal [759]) );
  inv U762 ( .a(n761), .out(\sig_prgm_register/or_signal [760]) );
  inv U763 ( .a(n762), .out(\sig_prgm_register/or_signal [761]) );
  inv U764 ( .a(n763), .out(\sig_prgm_register/or_signal [762]) );
  inv U765 ( .a(n764), .out(\sig_prgm_register/or_signal [763]) );
  inv U766 ( .a(n765), .out(\sig_prgm_register/or_signal [764]) );
  inv U767 ( .a(n766), .out(\sig_prgm_register/or_signal [765]) );
  inv U768 ( .a(n767), .out(\sig_prgm_register/or_signal [766]) );
  inv U769 ( .a(n768), .out(\sig_prgm_register/or_signal [767]) );
  inv U770 ( .a(n769), .out(\sig_prgm_register/or_signal [768]) );
  inv U771 ( .a(n770), .out(\sig_prgm_register/or_signal [769]) );
  inv U772 ( .a(n771), .out(\sig_prgm_register/or_signal [770]) );
  inv U773 ( .a(n772), .out(\sig_prgm_register/or_signal [771]) );
  inv U774 ( .a(n773), .out(\sig_prgm_register/or_signal [772]) );
  inv U775 ( .a(n774), .out(\sig_prgm_register/or_signal [773]) );
  inv U776 ( .a(n775), .out(\sig_prgm_register/or_signal [774]) );
  inv U777 ( .a(n776), .out(\sig_prgm_register/or_signal [775]) );
  inv U778 ( .a(n777), .out(\sig_prgm_register/or_signal [776]) );
  inv U779 ( .a(n778), .out(\sig_prgm_register/or_signal [777]) );
  inv U780 ( .a(n779), .out(\sig_prgm_register/or_signal [778]) );
  inv U781 ( .a(n780), .out(\sig_prgm_register/or_signal [779]) );
  inv U782 ( .a(n781), .out(\sig_prgm_register/or_signal [780]) );
  inv U783 ( .a(n782), .out(\sig_prgm_register/or_signal [781]) );
  inv U784 ( .a(n783), .out(\sig_prgm_register/or_signal [782]) );
  inv U785 ( .a(n784), .out(\sig_prgm_register/or_signal [783]) );
  inv U786 ( .a(n785), .out(\sig_prgm_register/or_signal [784]) );
  inv U787 ( .a(n786), .out(\sig_prgm_register/or_signal [785]) );
  inv U788 ( .a(n787), .out(\sig_prgm_register/or_signal [786]) );
  inv U789 ( .a(n788), .out(\sig_prgm_register/or_signal [787]) );
  inv U790 ( .a(n789), .out(\sig_prgm_register/or_signal [788]) );
  inv U791 ( .a(n790), .out(\sig_prgm_register/or_signal [789]) );
  inv U792 ( .a(n791), .out(\sig_prgm_register/or_signal [790]) );
  inv U793 ( .a(n792), .out(\sig_prgm_register/or_signal [791]) );
  inv U794 ( .a(n793), .out(\sig_prgm_register/or_signal [792]) );
  inv U795 ( .a(n794), .out(\sig_prgm_register/or_signal [793]) );
  inv U796 ( .a(n795), .out(\sig_prgm_register/or_signal [794]) );
  inv U797 ( .a(n796), .out(\sig_prgm_register/or_signal [795]) );
  inv U798 ( .a(n797), .out(\sig_prgm_register/or_signal [796]) );
  inv U799 ( .a(n798), .out(\sig_prgm_register/or_signal [797]) );
  inv U800 ( .a(n799), .out(\sig_prgm_register/or_signal [798]) );
  inv U801 ( .a(n800), .out(\sig_prgm_register/or_signal [799]) );
  inv U802 ( .a(n801), .out(\sig_prgm_register/or_signal [800]) );
  inv U803 ( .a(n802), .out(\sig_prgm_register/or_signal [801]) );
  inv U804 ( .a(n803), .out(\sig_prgm_register/or_signal [802]) );
  inv U805 ( .a(n804), .out(\sig_prgm_register/or_signal [803]) );
  inv U806 ( .a(n805), .out(\sig_prgm_register/or_signal [804]) );
  inv U807 ( .a(n806), .out(\sig_prgm_register/or_signal [805]) );
  inv U808 ( .a(n807), .out(\sig_prgm_register/or_signal [806]) );
  inv U809 ( .a(n808), .out(\sig_prgm_register/or_signal [807]) );
  inv U810 ( .a(n809), .out(\sig_prgm_register/or_signal [808]) );
  inv U811 ( .a(n810), .out(\sig_prgm_register/or_signal [809]) );
  inv U812 ( .a(n811), .out(\sig_prgm_register/or_signal [810]) );
  inv U813 ( .a(n812), .out(\sig_prgm_register/or_signal [811]) );
  inv U814 ( .a(n813), .out(\sig_prgm_register/or_signal [812]) );
  inv U815 ( .a(n814), .out(\sig_prgm_register/or_signal [813]) );
  inv U816 ( .a(n815), .out(\sig_prgm_register/or_signal [814]) );
  inv U817 ( .a(n816), .out(\sig_prgm_register/or_signal [815]) );
  inv U818 ( .a(n817), .out(\sig_prgm_register/or_signal [816]) );
  inv U819 ( .a(n818), .out(\sig_prgm_register/or_signal [817]) );
  inv U820 ( .a(n819), .out(\sig_prgm_register/or_signal [818]) );
  inv U821 ( .a(n820), .out(\sig_prgm_register/or_signal [819]) );
  inv U822 ( .a(n821), .out(\sig_prgm_register/or_signal [820]) );
  inv U823 ( .a(n822), .out(\sig_prgm_register/or_signal [821]) );
  inv U824 ( .a(n823), .out(\sig_prgm_register/or_signal [822]) );
  inv U825 ( .a(n824), .out(\sig_prgm_register/or_signal [823]) );
  inv U826 ( .a(n825), .out(\sig_prgm_register/or_signal [824]) );
  inv U827 ( .a(n826), .out(\sig_prgm_register/or_signal [825]) );
  inv U828 ( .a(n827), .out(\sig_prgm_register/or_signal [826]) );
  inv U829 ( .a(n828), .out(\sig_prgm_register/or_signal [827]) );
  inv U830 ( .a(n829), .out(\sig_prgm_register/or_signal [828]) );
  inv U831 ( .a(n830), .out(\sig_prgm_register/or_signal [829]) );
  inv U832 ( .a(n831), .out(\sig_prgm_register/or_signal [830]) );
  inv U833 ( .a(n832), .out(\sig_prgm_register/or_signal [831]) );
  inv U834 ( .a(n833), .out(\sig_prgm_register/or_signal [832]) );
  inv U835 ( .a(n834), .out(\sig_prgm_register/or_signal [833]) );
  inv U836 ( .a(n835), .out(\sig_prgm_register/or_signal [834]) );
  inv U837 ( .a(n836), .out(\sig_prgm_register/or_signal [835]) );
  inv U838 ( .a(n837), .out(\sig_prgm_register/or_signal [836]) );
  inv U839 ( .a(n838), .out(\sig_prgm_register/or_signal [837]) );
  inv U840 ( .a(n839), .out(\sig_prgm_register/or_signal [838]) );
  inv U841 ( .a(n840), .out(\sig_prgm_register/or_signal [839]) );
  inv U842 ( .a(n841), .out(\sig_prgm_register/or_signal [840]) );
  inv U843 ( .a(n842), .out(\sig_prgm_register/or_signal [841]) );
  inv U844 ( .a(n843), .out(\sig_prgm_register/or_signal [842]) );
  inv U845 ( .a(n844), .out(\sig_prgm_register/or_signal [843]) );
  inv U846 ( .a(n845), .out(\sig_prgm_register/or_signal [844]) );
  inv U847 ( .a(n846), .out(\sig_prgm_register/or_signal [845]) );
  inv U848 ( .a(n847), .out(\sig_prgm_register/or_signal [846]) );
  inv U849 ( .a(n848), .out(\sig_prgm_register/or_signal [847]) );
  inv U850 ( .a(n849), .out(\sig_prgm_register/or_signal [848]) );
  inv U851 ( .a(n850), .out(\sig_prgm_register/or_signal [849]) );
  inv U852 ( .a(n851), .out(\sig_prgm_register/or_signal [850]) );
  inv U853 ( .a(n852), .out(\sig_prgm_register/or_signal [851]) );
  inv U854 ( .a(n853), .out(\sig_prgm_register/or_signal [852]) );
  inv U855 ( .a(n854), .out(\sig_prgm_register/or_signal [853]) );
  inv U856 ( .a(n855), .out(\sig_prgm_register/or_signal [854]) );
  inv U857 ( .a(n856), .out(\sig_prgm_register/or_signal [855]) );
  inv U858 ( .a(n857), .out(\sig_prgm_register/or_signal [856]) );
  inv U859 ( .a(n858), .out(\sig_prgm_register/or_signal [857]) );
  inv U860 ( .a(n859), .out(\sig_prgm_register/or_signal [858]) );
  inv U861 ( .a(n860), .out(\sig_prgm_register/or_signal [859]) );
  inv U862 ( .a(n861), .out(\sig_prgm_register/or_signal [860]) );
  inv U863 ( .a(n862), .out(\sig_prgm_register/or_signal [861]) );
  inv U864 ( .a(n863), .out(\sig_prgm_register/or_signal [862]) );
  inv U865 ( .a(n864), .out(\sig_prgm_register/or_signal [863]) );
  inv U866 ( .a(n865), .out(\sig_prgm_register/or_signal [864]) );
  inv U867 ( .a(n866), .out(\sig_prgm_register/or_signal [865]) );
  inv U868 ( .a(n867), .out(\sig_prgm_register/or_signal [866]) );
  inv U869 ( .a(n868), .out(\sig_prgm_register/or_signal [867]) );
  inv U870 ( .a(n869), .out(\sig_prgm_register/or_signal [868]) );
  inv U871 ( .a(n870), .out(\sig_prgm_register/or_signal [869]) );
  inv U872 ( .a(n871), .out(\sig_prgm_register/or_signal [870]) );
  inv U873 ( .a(n872), .out(\sig_prgm_register/or_signal [871]) );
  inv U874 ( .a(n873), .out(\sig_prgm_register/or_signal [872]) );
  inv U875 ( .a(n874), .out(\sig_prgm_register/or_signal [873]) );
  inv U876 ( .a(n875), .out(\sig_prgm_register/or_signal [874]) );
  inv U877 ( .a(n876), .out(\sig_prgm_register/or_signal [875]) );
  inv U878 ( .a(n877), .out(\sig_prgm_register/or_signal [876]) );
  inv U879 ( .a(n878), .out(\sig_prgm_register/or_signal [877]) );
  inv U880 ( .a(n879), .out(\sig_prgm_register/or_signal [878]) );
  inv U881 ( .a(n880), .out(\sig_prgm_register/or_signal [879]) );
  inv U882 ( .a(n881), .out(\sig_prgm_register/or_signal [880]) );
  inv U883 ( .a(n882), .out(\sig_prgm_register/or_signal [881]) );
  inv U884 ( .a(n883), .out(\sig_prgm_register/or_signal [882]) );
  inv U885 ( .a(n884), .out(\sig_prgm_register/or_signal [883]) );
  inv U886 ( .a(n885), .out(\sig_prgm_register/or_signal [884]) );
  inv U887 ( .a(n886), .out(\sig_prgm_register/or_signal [885]) );
  inv U888 ( .a(n887), .out(\sig_prgm_register/or_signal [886]) );
  inv U889 ( .a(n888), .out(\sig_prgm_register/or_signal [887]) );
  inv U890 ( .a(n889), .out(\sig_prgm_register/or_signal [888]) );
  inv U891 ( .a(n890), .out(\sig_prgm_register/or_signal [889]) );
  inv U892 ( .a(n891), .out(\sig_prgm_register/or_signal [890]) );
  inv U893 ( .a(n892), .out(\sig_prgm_register/or_signal [891]) );
  inv U894 ( .a(n893), .out(\sig_prgm_register/or_signal [892]) );
  inv U895 ( .a(n894), .out(\sig_prgm_register/or_signal [893]) );
  inv U896 ( .a(n895), .out(\sig_prgm_register/or_signal [894]) );
  inv U897 ( .a(n896), .out(\sig_prgm_register/or_signal [895]) );
  inv U898 ( .a(n897), .out(\sig_prgm_register/or_signal [896]) );
  inv U899 ( .a(n898), .out(\sig_prgm_register/or_signal [897]) );
  inv U900 ( .a(n899), .out(\sig_prgm_register/or_signal [898]) );
  inv U901 ( .a(n900), .out(\sig_prgm_register/or_signal [899]) );
  inv U902 ( .a(n901), .out(\sig_prgm_register/or_signal [900]) );
  inv U903 ( .a(n902), .out(\sig_prgm_register/or_signal [901]) );
  inv U904 ( .a(n903), .out(\sig_prgm_register/or_signal [902]) );
  inv U905 ( .a(n904), .out(\sig_prgm_register/or_signal [903]) );
  inv U906 ( .a(n905), .out(\sig_prgm_register/or_signal [904]) );
  inv U907 ( .a(n906), .out(\sig_prgm_register/or_signal [905]) );
  inv U908 ( .a(n907), .out(\sig_prgm_register/or_signal [906]) );
  inv U909 ( .a(n908), .out(\sig_prgm_register/or_signal [907]) );
  inv U910 ( .a(n909), .out(\sig_prgm_register/or_signal [908]) );
  inv U911 ( .a(n910), .out(\sig_prgm_register/or_signal [909]) );
  inv U912 ( .a(n911), .out(\sig_prgm_register/or_signal [910]) );
  inv U913 ( .a(n912), .out(\sig_prgm_register/or_signal [911]) );
  inv U914 ( .a(n913), .out(\sig_prgm_register/or_signal [912]) );
  inv U915 ( .a(n914), .out(\sig_prgm_register/or_signal [913]) );
  inv U916 ( .a(n915), .out(\sig_prgm_register/or_signal [914]) );
  inv U917 ( .a(n916), .out(\sig_prgm_register/or_signal [915]) );
  inv U918 ( .a(n917), .out(\sig_prgm_register/or_signal [916]) );
  inv U919 ( .a(n918), .out(\sig_prgm_register/or_signal [917]) );
  inv U920 ( .a(n919), .out(\sig_prgm_register/or_signal [918]) );
  inv U921 ( .a(n920), .out(\sig_prgm_register/or_signal [919]) );
  inv U922 ( .a(n921), .out(\sig_prgm_register/or_signal [920]) );
  inv U923 ( .a(n922), .out(\sig_prgm_register/or_signal [921]) );
  inv U924 ( .a(n923), .out(\sig_prgm_register/or_signal [922]) );
  inv U925 ( .a(n924), .out(\sig_prgm_register/or_signal [923]) );
  inv U926 ( .a(n925), .out(\sig_prgm_register/or_signal [924]) );
  inv U927 ( .a(n926), .out(\sig_prgm_register/or_signal [925]) );
  inv U928 ( .a(n927), .out(\sig_prgm_register/or_signal [926]) );
  inv U929 ( .a(n928), .out(\sig_prgm_register/or_signal [927]) );
  inv U930 ( .a(n929), .out(\sig_prgm_register/or_signal [928]) );
  inv U931 ( .a(n930), .out(\sig_prgm_register/or_signal [929]) );
  inv U932 ( .a(n931), .out(\sig_prgm_register/or_signal [930]) );
  inv U933 ( .a(n932), .out(\sig_prgm_register/or_signal [931]) );
  inv U934 ( .a(n933), .out(\sig_prgm_register/or_signal [932]) );
  inv U935 ( .a(n934), .out(\sig_prgm_register/or_signal [933]) );
  inv U936 ( .a(n935), .out(\sig_prgm_register/or_signal [934]) );
  inv U937 ( .a(n936), .out(\sig_prgm_register/or_signal [935]) );
  inv U938 ( .a(n937), .out(\sig_prgm_register/or_signal [936]) );
  inv U939 ( .a(n938), .out(\sig_prgm_register/or_signal [937]) );
  inv U940 ( .a(n939), .out(\sig_prgm_register/or_signal [938]) );
  inv U941 ( .a(n940), .out(\sig_prgm_register/or_signal [939]) );
  inv U942 ( .a(n941), .out(\sig_prgm_register/or_signal [940]) );
  inv U943 ( .a(n942), .out(\sig_prgm_register/or_signal [941]) );
  inv U944 ( .a(n943), .out(\sig_prgm_register/or_signal [942]) );
  inv U945 ( .a(n944), .out(\sig_prgm_register/or_signal [943]) );
  inv U946 ( .a(n945), .out(\sig_prgm_register/or_signal [944]) );
  inv U947 ( .a(n946), .out(\sig_prgm_register/or_signal [945]) );
  inv U948 ( .a(n947), .out(\sig_prgm_register/or_signal [946]) );
  inv U949 ( .a(n948), .out(\sig_prgm_register/or_signal [947]) );
  inv U950 ( .a(n949), .out(\sig_prgm_register/or_signal [948]) );
  inv U951 ( .a(n950), .out(\sig_prgm_register/or_signal [949]) );
  inv U952 ( .a(n951), .out(\sig_prgm_register/or_signal [950]) );
  inv U953 ( .a(n952), .out(\sig_prgm_register/or_signal [951]) );
  inv U954 ( .a(n953), .out(\sig_prgm_register/or_signal [952]) );
  inv U955 ( .a(n954), .out(\sig_prgm_register/or_signal [953]) );
  inv U956 ( .a(n955), .out(\sig_prgm_register/or_signal [954]) );
  inv U957 ( .a(n956), .out(\sig_prgm_register/or_signal [955]) );
  inv U958 ( .a(n957), .out(\sig_prgm_register/or_signal [956]) );
  inv U959 ( .a(n958), .out(\sig_prgm_register/or_signal [957]) );
  inv U960 ( .a(n959), .out(\sig_prgm_register/or_signal [958]) );
  inv U961 ( .a(n960), .out(\sig_prgm_register/or_signal [959]) );
  inv U962 ( .a(n961), .out(\sig_prgm_register/or_signal [960]) );
  inv U963 ( .a(n962), .out(\sig_prgm_register/or_signal [961]) );
  inv U964 ( .a(n963), .out(\sig_prgm_register/or_signal [962]) );
  inv U965 ( .a(n964), .out(\sig_prgm_register/or_signal [963]) );
  inv U966 ( .a(n965), .out(\sig_prgm_register/or_signal [964]) );
  inv U967 ( .a(n966), .out(\sig_prgm_register/or_signal [965]) );
  inv U968 ( .a(n967), .out(\sig_prgm_register/or_signal [966]) );
  inv U969 ( .a(n968), .out(\sig_prgm_register/or_signal [967]) );
  inv U970 ( .a(n969), .out(\sig_prgm_register/or_signal [968]) );
  inv U971 ( .a(n970), .out(\sig_prgm_register/or_signal [969]) );
  inv U972 ( .a(n971), .out(\sig_prgm_register/or_signal [970]) );
  inv U973 ( .a(n972), .out(\sig_prgm_register/or_signal [971]) );
  inv U974 ( .a(n973), .out(\sig_prgm_register/or_signal [972]) );
  inv U975 ( .a(n974), .out(\sig_prgm_register/or_signal [973]) );
  inv U976 ( .a(n975), .out(\sig_prgm_register/or_signal [974]) );
  inv U977 ( .a(n976), .out(\sig_prgm_register/or_signal [975]) );
  inv U978 ( .a(n977), .out(\sig_prgm_register/or_signal [976]) );
  inv U979 ( .a(n978), .out(\sig_prgm_register/or_signal [977]) );
  inv U980 ( .a(n979), .out(\sig_prgm_register/or_signal [978]) );
  inv U981 ( .a(n980), .out(\sig_prgm_register/or_signal [979]) );
  inv U982 ( .a(n981), .out(\sig_prgm_register/or_signal [980]) );
  inv U983 ( .a(n982), .out(\sig_prgm_register/or_signal [981]) );
  inv U984 ( .a(n983), .out(\sig_prgm_register/or_signal [982]) );
  inv U985 ( .a(n984), .out(\sig_prgm_register/or_signal [983]) );
  inv U986 ( .a(n985), .out(\sig_prgm_register/or_signal [984]) );
  inv U987 ( .a(n986), .out(\sig_prgm_register/or_signal [985]) );
  inv U988 ( .a(n987), .out(\sig_prgm_register/or_signal [986]) );
  inv U989 ( .a(n988), .out(\sig_prgm_register/or_signal [987]) );
  inv U990 ( .a(n989), .out(\sig_prgm_register/or_signal [988]) );
  inv U991 ( .a(n990), .out(\sig_prgm_register/or_signal [989]) );
  inv U992 ( .a(n991), .out(\sig_prgm_register/or_signal [990]) );
  inv U993 ( .a(n992), .out(\sig_prgm_register/or_signal [991]) );
  inv U994 ( .a(n993), .out(\sig_prgm_register/or_signal [992]) );
  inv U995 ( .a(n994), .out(\sig_prgm_register/or_signal [993]) );
  inv U996 ( .a(n995), .out(\sig_prgm_register/or_signal [994]) );
  inv U997 ( .a(n996), .out(\sig_prgm_register/or_signal [995]) );
  inv U998 ( .a(n997), .out(\sig_prgm_register/or_signal [996]) );
  inv U999 ( .a(n998), .out(\sig_prgm_register/or_signal [997]) );
  inv U1000 ( .a(n999), .out(\sig_prgm_register/or_signal [998]) );
  inv U1001 ( .a(n1000), .out(\sig_prgm_register/or_signal [999]) );
  inv U1002 ( .a(n1001), .out(\sig_prgm_register/or_signal [1000]) );
  inv U1003 ( .a(n1002), .out(\sig_prgm_register/or_signal [1001]) );
  inv U1004 ( .a(n1003), .out(\sig_prgm_register/or_signal [1002]) );
  inv U1005 ( .a(n1004), .out(\sig_prgm_register/or_signal [1003]) );
  inv U1006 ( .a(n1005), .out(\sig_prgm_register/or_signal [1004]) );
  inv U1007 ( .a(n1006), .out(\sig_prgm_register/or_signal [1005]) );
  inv U1008 ( .a(n1007), .out(\sig_prgm_register/or_signal [1006]) );
  inv U1009 ( .a(n1008), .out(\sig_prgm_register/or_signal [1007]) );
  inv U1010 ( .a(n1009), .out(\sig_prgm_register/or_signal [1008]) );
  inv U1011 ( .a(n1010), .out(\sig_prgm_register/or_signal [1009]) );
  inv U1012 ( .a(n1011), .out(\sig_prgm_register/or_signal [1010]) );
  inv U1013 ( .a(n1012), .out(\sig_prgm_register/or_signal [1011]) );
  inv U1014 ( .a(n1013), .out(\sig_prgm_register/or_signal [1012]) );
  inv U1015 ( .a(n1014), .out(\sig_prgm_register/or_signal [1013]) );
  inv U1016 ( .a(n1015), .out(\sig_prgm_register/or_signal [1014]) );
  inv U1017 ( .a(n1016), .out(\sig_prgm_register/or_signal [1015]) );
  inv U1018 ( .a(n1017), .out(\sig_prgm_register/or_signal [1016]) );
  inv U1019 ( .a(n1018), .out(\sig_prgm_register/or_signal [1017]) );
  inv U1020 ( .a(n1019), .out(\sig_prgm_register/or_signal [1018]) );
  inv U1021 ( .a(n1020), .out(\sig_prgm_register/or_signal [1019]) );
  inv U1022 ( .a(n1021), .out(\sig_prgm_register/or_signal [1020]) );
  inv U1023 ( .a(n1022), .out(\sig_prgm_register/or_signal [1021]) );
  inv U1024 ( .a(n1023), .out(\sig_prgm_register/or_signal [1022]) );
  inv U1025 ( .a(n1024), .out(\sig_prgm_register/or_signal [1023]) );
  inv U1026 ( .a(sig), .out(n1) );
  inv U1027 ( .a(b[0]), .out(n2) );
  inv U1028 ( .a(b[1]), .out(n3) );
  inv U1029 ( .a(b[2]), .out(n4) );
  inv U1030 ( .a(b[3]), .out(n5) );
  inv U1031 ( .a(b[4]), .out(n6) );
  inv U1032 ( .a(b[5]), .out(n7) );
  inv U1033 ( .a(b[6]), .out(n8) );
  inv U1034 ( .a(b[7]), .out(n9) );
  inv U1035 ( .a(b[8]), .out(n10) );
  inv U1036 ( .a(b[9]), .out(n11) );
  inv U1037 ( .a(b[10]), .out(n12) );
  inv U1038 ( .a(b[11]), .out(n13) );
  inv U1039 ( .a(b[12]), .out(n14) );
  inv U1040 ( .a(b[13]), .out(n15) );
  inv U1041 ( .a(b[14]), .out(n16) );
  inv U1042 ( .a(b[15]), .out(n17) );
  inv U1043 ( .a(b[16]), .out(n18) );
  inv U1044 ( .a(b[17]), .out(n19) );
  inv U1045 ( .a(b[18]), .out(n20) );
  inv U1046 ( .a(b[19]), .out(n21) );
  inv U1047 ( .a(b[20]), .out(n22) );
  inv U1048 ( .a(b[21]), .out(n23) );
  inv U1049 ( .a(b[22]), .out(n24) );
  inv U1050 ( .a(b[23]), .out(n25) );
  inv U1051 ( .a(b[24]), .out(n26) );
  inv U1052 ( .a(b[25]), .out(n27) );
  inv U1053 ( .a(b[26]), .out(n28) );
  inv U1054 ( .a(b[27]), .out(n29) );
  inv U1055 ( .a(b[28]), .out(n30) );
  inv U1056 ( .a(b[29]), .out(n31) );
  inv U1057 ( .a(b[30]), .out(n32) );
  inv U1058 ( .a(b[31]), .out(n33) );
  inv U1059 ( .a(b[32]), .out(n34) );
  inv U1060 ( .a(b[33]), .out(n35) );
  inv U1061 ( .a(b[34]), .out(n36) );
  inv U1062 ( .a(b[35]), .out(n37) );
  inv U1063 ( .a(b[36]), .out(n38) );
  inv U1064 ( .a(b[37]), .out(n39) );
  inv U1065 ( .a(b[38]), .out(n40) );
  inv U1066 ( .a(b[39]), .out(n41) );
  inv U1067 ( .a(b[40]), .out(n42) );
  inv U1068 ( .a(b[41]), .out(n43) );
  inv U1069 ( .a(b[42]), .out(n44) );
  inv U1070 ( .a(b[43]), .out(n45) );
  inv U1071 ( .a(b[44]), .out(n46) );
  inv U1072 ( .a(b[45]), .out(n47) );
  inv U1073 ( .a(b[46]), .out(n48) );
  inv U1074 ( .a(b[47]), .out(n49) );
  inv U1075 ( .a(b[48]), .out(n50) );
  inv U1076 ( .a(b[49]), .out(n51) );
  inv U1077 ( .a(b[50]), .out(n52) );
  inv U1078 ( .a(b[51]), .out(n53) );
  inv U1079 ( .a(b[52]), .out(n54) );
  inv U1080 ( .a(b[53]), .out(n55) );
  inv U1081 ( .a(b[54]), .out(n56) );
  inv U1082 ( .a(b[55]), .out(n57) );
  inv U1083 ( .a(b[56]), .out(n58) );
  inv U1084 ( .a(b[57]), .out(n59) );
  inv U1085 ( .a(b[58]), .out(n60) );
  inv U1086 ( .a(b[59]), .out(n61) );
  inv U1087 ( .a(b[60]), .out(n62) );
  inv U1088 ( .a(b[61]), .out(n63) );
  inv U1089 ( .a(b[62]), .out(n64) );
  inv U1090 ( .a(b[63]), .out(n65) );
  inv U1091 ( .a(b[64]), .out(n66) );
  inv U1092 ( .a(b[65]), .out(n67) );
  inv U1093 ( .a(b[66]), .out(n68) );
  inv U1094 ( .a(b[67]), .out(n69) );
  inv U1095 ( .a(b[68]), .out(n70) );
  inv U1096 ( .a(b[69]), .out(n71) );
  inv U1097 ( .a(b[70]), .out(n72) );
  inv U1098 ( .a(b[71]), .out(n73) );
  inv U1099 ( .a(b[72]), .out(n74) );
  inv U1100 ( .a(b[73]), .out(n75) );
  inv U1101 ( .a(b[74]), .out(n76) );
  inv U1102 ( .a(b[75]), .out(n77) );
  inv U1103 ( .a(b[76]), .out(n78) );
  inv U1104 ( .a(b[77]), .out(n79) );
  inv U1105 ( .a(b[78]), .out(n80) );
  inv U1106 ( .a(b[79]), .out(n81) );
  inv U1107 ( .a(b[80]), .out(n82) );
  inv U1108 ( .a(b[81]), .out(n83) );
  inv U1109 ( .a(b[82]), .out(n84) );
  inv U1110 ( .a(b[83]), .out(n85) );
  inv U1111 ( .a(b[84]), .out(n86) );
  inv U1112 ( .a(b[85]), .out(n87) );
  inv U1113 ( .a(b[86]), .out(n88) );
  inv U1114 ( .a(b[87]), .out(n89) );
  inv U1115 ( .a(b[88]), .out(n90) );
  inv U1116 ( .a(b[89]), .out(n91) );
  inv U1117 ( .a(b[90]), .out(n92) );
  inv U1118 ( .a(b[91]), .out(n93) );
  inv U1119 ( .a(b[92]), .out(n94) );
  inv U1120 ( .a(b[93]), .out(n95) );
  inv U1121 ( .a(b[94]), .out(n96) );
  inv U1122 ( .a(b[95]), .out(n97) );
  inv U1123 ( .a(b[96]), .out(n98) );
  inv U1124 ( .a(b[97]), .out(n99) );
  inv U1125 ( .a(b[98]), .out(n100) );
  inv U1126 ( .a(b[99]), .out(n101) );
  inv U1127 ( .a(b[100]), .out(n102) );
  inv U1128 ( .a(b[101]), .out(n103) );
  inv U1129 ( .a(b[102]), .out(n104) );
  inv U1130 ( .a(b[103]), .out(n105) );
  inv U1131 ( .a(b[104]), .out(n106) );
  inv U1132 ( .a(b[105]), .out(n107) );
  inv U1133 ( .a(b[106]), .out(n108) );
  inv U1134 ( .a(b[107]), .out(n109) );
  inv U1135 ( .a(b[108]), .out(n110) );
  inv U1136 ( .a(b[109]), .out(n111) );
  inv U1137 ( .a(b[110]), .out(n112) );
  inv U1138 ( .a(b[111]), .out(n113) );
  inv U1139 ( .a(b[112]), .out(n114) );
  inv U1140 ( .a(b[113]), .out(n115) );
  inv U1141 ( .a(b[114]), .out(n116) );
  inv U1142 ( .a(b[115]), .out(n117) );
  inv U1143 ( .a(b[116]), .out(n118) );
  inv U1144 ( .a(b[117]), .out(n119) );
  inv U1145 ( .a(b[118]), .out(n120) );
  inv U1146 ( .a(b[119]), .out(n121) );
  inv U1147 ( .a(b[120]), .out(n122) );
  inv U1148 ( .a(b[121]), .out(n123) );
  inv U1149 ( .a(b[122]), .out(n124) );
  inv U1150 ( .a(b[123]), .out(n125) );
  inv U1151 ( .a(b[124]), .out(n126) );
  inv U1152 ( .a(b[125]), .out(n127) );
  inv U1153 ( .a(b[126]), .out(n128) );
  inv U1154 ( .a(b[127]), .out(n129) );
  inv U1155 ( .a(b[128]), .out(n130) );
  inv U1156 ( .a(b[129]), .out(n131) );
  inv U1157 ( .a(b[130]), .out(n132) );
  inv U1158 ( .a(b[131]), .out(n133) );
  inv U1159 ( .a(b[132]), .out(n134) );
  inv U1160 ( .a(b[133]), .out(n135) );
  inv U1161 ( .a(b[134]), .out(n136) );
  inv U1162 ( .a(b[135]), .out(n137) );
  inv U1163 ( .a(b[136]), .out(n138) );
  inv U1164 ( .a(b[137]), .out(n139) );
  inv U1165 ( .a(b[138]), .out(n140) );
  inv U1166 ( .a(b[139]), .out(n141) );
  inv U1167 ( .a(b[140]), .out(n142) );
  inv U1168 ( .a(b[141]), .out(n143) );
  inv U1169 ( .a(b[142]), .out(n144) );
  inv U1170 ( .a(b[143]), .out(n145) );
  inv U1171 ( .a(b[144]), .out(n146) );
  inv U1172 ( .a(b[145]), .out(n147) );
  inv U1173 ( .a(b[146]), .out(n148) );
  inv U1174 ( .a(b[147]), .out(n149) );
  inv U1175 ( .a(b[148]), .out(n150) );
  inv U1176 ( .a(b[149]), .out(n151) );
  inv U1177 ( .a(b[150]), .out(n152) );
  inv U1178 ( .a(b[151]), .out(n153) );
  inv U1179 ( .a(b[152]), .out(n154) );
  inv U1180 ( .a(b[153]), .out(n155) );
  inv U1181 ( .a(b[154]), .out(n156) );
  inv U1182 ( .a(b[155]), .out(n157) );
  inv U1183 ( .a(b[156]), .out(n158) );
  inv U1184 ( .a(b[157]), .out(n159) );
  inv U1185 ( .a(b[158]), .out(n160) );
  inv U1186 ( .a(b[159]), .out(n161) );
  inv U1187 ( .a(b[160]), .out(n162) );
  inv U1188 ( .a(b[161]), .out(n163) );
  inv U1189 ( .a(b[162]), .out(n164) );
  inv U1190 ( .a(b[163]), .out(n165) );
  inv U1191 ( .a(b[164]), .out(n166) );
  inv U1192 ( .a(b[165]), .out(n167) );
  inv U1193 ( .a(b[166]), .out(n168) );
  inv U1194 ( .a(b[167]), .out(n169) );
  inv U1195 ( .a(b[168]), .out(n170) );
  inv U1196 ( .a(b[169]), .out(n171) );
  inv U1197 ( .a(b[170]), .out(n172) );
  inv U1198 ( .a(b[171]), .out(n173) );
  inv U1199 ( .a(b[172]), .out(n174) );
  inv U1200 ( .a(b[173]), .out(n175) );
  inv U1201 ( .a(b[174]), .out(n176) );
  inv U1202 ( .a(b[175]), .out(n177) );
  inv U1203 ( .a(b[176]), .out(n178) );
  inv U1204 ( .a(b[177]), .out(n179) );
  inv U1205 ( .a(b[178]), .out(n180) );
  inv U1206 ( .a(b[179]), .out(n181) );
  inv U1207 ( .a(b[180]), .out(n182) );
  inv U1208 ( .a(b[181]), .out(n183) );
  inv U1209 ( .a(b[182]), .out(n184) );
  inv U1210 ( .a(b[183]), .out(n185) );
  inv U1211 ( .a(b[184]), .out(n186) );
  inv U1212 ( .a(b[185]), .out(n187) );
  inv U1213 ( .a(b[186]), .out(n188) );
  inv U1214 ( .a(b[187]), .out(n189) );
  inv U1215 ( .a(b[188]), .out(n190) );
  inv U1216 ( .a(b[189]), .out(n191) );
  inv U1217 ( .a(b[190]), .out(n192) );
  inv U1218 ( .a(b[191]), .out(n193) );
  inv U1219 ( .a(b[192]), .out(n194) );
  inv U1220 ( .a(b[193]), .out(n195) );
  inv U1221 ( .a(b[194]), .out(n196) );
  inv U1222 ( .a(b[195]), .out(n197) );
  inv U1223 ( .a(b[196]), .out(n198) );
  inv U1224 ( .a(b[197]), .out(n199) );
  inv U1225 ( .a(b[198]), .out(n200) );
  inv U1226 ( .a(b[199]), .out(n201) );
  inv U1227 ( .a(b[200]), .out(n202) );
  inv U1228 ( .a(b[201]), .out(n203) );
  inv U1229 ( .a(b[202]), .out(n204) );
  inv U1230 ( .a(b[203]), .out(n205) );
  inv U1231 ( .a(b[204]), .out(n206) );
  inv U1232 ( .a(b[205]), .out(n207) );
  inv U1233 ( .a(b[206]), .out(n208) );
  inv U1234 ( .a(b[207]), .out(n209) );
  inv U1235 ( .a(b[208]), .out(n210) );
  inv U1236 ( .a(b[209]), .out(n211) );
  inv U1237 ( .a(b[210]), .out(n212) );
  inv U1238 ( .a(b[211]), .out(n213) );
  inv U1239 ( .a(b[212]), .out(n214) );
  inv U1240 ( .a(b[213]), .out(n215) );
  inv U1241 ( .a(b[214]), .out(n216) );
  inv U1242 ( .a(b[215]), .out(n217) );
  inv U1243 ( .a(b[216]), .out(n218) );
  inv U1244 ( .a(b[217]), .out(n219) );
  inv U1245 ( .a(b[218]), .out(n220) );
  inv U1246 ( .a(b[219]), .out(n221) );
  inv U1247 ( .a(b[220]), .out(n222) );
  inv U1248 ( .a(b[221]), .out(n223) );
  inv U1249 ( .a(b[222]), .out(n224) );
  inv U1250 ( .a(b[223]), .out(n225) );
  inv U1251 ( .a(b[224]), .out(n226) );
  inv U1252 ( .a(b[225]), .out(n227) );
  inv U1253 ( .a(b[226]), .out(n228) );
  inv U1254 ( .a(b[227]), .out(n229) );
  inv U1255 ( .a(b[228]), .out(n230) );
  inv U1256 ( .a(b[229]), .out(n231) );
  inv U1257 ( .a(b[230]), .out(n232) );
  inv U1258 ( .a(b[231]), .out(n233) );
  inv U1259 ( .a(b[232]), .out(n234) );
  inv U1260 ( .a(b[233]), .out(n235) );
  inv U1261 ( .a(b[234]), .out(n236) );
  inv U1262 ( .a(b[235]), .out(n237) );
  inv U1263 ( .a(b[236]), .out(n238) );
  inv U1264 ( .a(b[237]), .out(n239) );
  inv U1265 ( .a(b[238]), .out(n240) );
  inv U1266 ( .a(b[239]), .out(n241) );
  inv U1267 ( .a(b[240]), .out(n242) );
  inv U1268 ( .a(b[241]), .out(n243) );
  inv U1269 ( .a(b[242]), .out(n244) );
  inv U1270 ( .a(b[243]), .out(n245) );
  inv U1271 ( .a(b[244]), .out(n246) );
  inv U1272 ( .a(b[245]), .out(n247) );
  inv U1273 ( .a(b[246]), .out(n248) );
  inv U1274 ( .a(b[247]), .out(n249) );
  inv U1275 ( .a(b[248]), .out(n250) );
  inv U1276 ( .a(b[249]), .out(n251) );
  inv U1277 ( .a(b[250]), .out(n252) );
  inv U1278 ( .a(b[251]), .out(n253) );
  inv U1279 ( .a(b[252]), .out(n254) );
  inv U1280 ( .a(b[253]), .out(n255) );
  inv U1281 ( .a(b[254]), .out(n256) );
  inv U1282 ( .a(b[255]), .out(n257) );
  inv U1283 ( .a(b[256]), .out(n258) );
  inv U1284 ( .a(b[257]), .out(n259) );
  inv U1285 ( .a(b[258]), .out(n260) );
  inv U1286 ( .a(b[259]), .out(n261) );
  inv U1287 ( .a(b[260]), .out(n262) );
  inv U1288 ( .a(b[261]), .out(n263) );
  inv U1289 ( .a(b[262]), .out(n264) );
  inv U1290 ( .a(b[263]), .out(n265) );
  inv U1291 ( .a(b[264]), .out(n266) );
  inv U1292 ( .a(b[265]), .out(n267) );
  inv U1293 ( .a(b[266]), .out(n268) );
  inv U1294 ( .a(b[267]), .out(n269) );
  inv U1295 ( .a(b[268]), .out(n270) );
  inv U1296 ( .a(b[269]), .out(n271) );
  inv U1297 ( .a(b[270]), .out(n272) );
  inv U1298 ( .a(b[271]), .out(n273) );
  inv U1299 ( .a(b[272]), .out(n274) );
  inv U1300 ( .a(b[273]), .out(n275) );
  inv U1301 ( .a(b[274]), .out(n276) );
  inv U1302 ( .a(b[275]), .out(n277) );
  inv U1303 ( .a(b[276]), .out(n278) );
  inv U1304 ( .a(b[277]), .out(n279) );
  inv U1305 ( .a(b[278]), .out(n280) );
  inv U1306 ( .a(b[279]), .out(n281) );
  inv U1307 ( .a(b[280]), .out(n282) );
  inv U1308 ( .a(b[281]), .out(n283) );
  inv U1309 ( .a(b[282]), .out(n284) );
  inv U1310 ( .a(b[283]), .out(n285) );
  inv U1311 ( .a(b[284]), .out(n286) );
  inv U1312 ( .a(b[285]), .out(n287) );
  inv U1313 ( .a(b[286]), .out(n288) );
  inv U1314 ( .a(b[287]), .out(n289) );
  inv U1315 ( .a(b[288]), .out(n290) );
  inv U1316 ( .a(b[289]), .out(n291) );
  inv U1317 ( .a(b[290]), .out(n292) );
  inv U1318 ( .a(b[291]), .out(n293) );
  inv U1319 ( .a(b[292]), .out(n294) );
  inv U1320 ( .a(b[293]), .out(n295) );
  inv U1321 ( .a(b[294]), .out(n296) );
  inv U1322 ( .a(b[295]), .out(n297) );
  inv U1323 ( .a(b[296]), .out(n298) );
  inv U1324 ( .a(b[297]), .out(n299) );
  inv U1325 ( .a(b[298]), .out(n300) );
  inv U1326 ( .a(b[299]), .out(n301) );
  inv U1327 ( .a(b[300]), .out(n302) );
  inv U1328 ( .a(b[301]), .out(n303) );
  inv U1329 ( .a(b[302]), .out(n304) );
  inv U1330 ( .a(b[303]), .out(n305) );
  inv U1331 ( .a(b[304]), .out(n306) );
  inv U1332 ( .a(b[305]), .out(n307) );
  inv U1333 ( .a(b[306]), .out(n308) );
  inv U1334 ( .a(b[307]), .out(n309) );
  inv U1335 ( .a(b[308]), .out(n310) );
  inv U1336 ( .a(b[309]), .out(n311) );
  inv U1337 ( .a(b[310]), .out(n312) );
  inv U1338 ( .a(b[311]), .out(n313) );
  inv U1339 ( .a(b[312]), .out(n314) );
  inv U1340 ( .a(b[313]), .out(n315) );
  inv U1341 ( .a(b[314]), .out(n316) );
  inv U1342 ( .a(b[315]), .out(n317) );
  inv U1343 ( .a(b[316]), .out(n318) );
  inv U1344 ( .a(b[317]), .out(n319) );
  inv U1345 ( .a(b[318]), .out(n320) );
  inv U1346 ( .a(b[319]), .out(n321) );
  inv U1347 ( .a(b[320]), .out(n322) );
  inv U1348 ( .a(b[321]), .out(n323) );
  inv U1349 ( .a(b[322]), .out(n324) );
  inv U1350 ( .a(b[323]), .out(n325) );
  inv U1351 ( .a(b[324]), .out(n326) );
  inv U1352 ( .a(b[325]), .out(n327) );
  inv U1353 ( .a(b[326]), .out(n328) );
  inv U1354 ( .a(b[327]), .out(n329) );
  inv U1355 ( .a(b[328]), .out(n330) );
  inv U1356 ( .a(b[329]), .out(n331) );
  inv U1357 ( .a(b[330]), .out(n332) );
  inv U1358 ( .a(b[331]), .out(n333) );
  inv U1359 ( .a(b[332]), .out(n334) );
  inv U1360 ( .a(b[333]), .out(n335) );
  inv U1361 ( .a(b[334]), .out(n336) );
  inv U1362 ( .a(b[335]), .out(n337) );
  inv U1363 ( .a(b[336]), .out(n338) );
  inv U1364 ( .a(b[337]), .out(n339) );
  inv U1365 ( .a(b[338]), .out(n340) );
  inv U1366 ( .a(b[339]), .out(n341) );
  inv U1367 ( .a(b[340]), .out(n342) );
  inv U1368 ( .a(b[341]), .out(n343) );
  inv U1369 ( .a(b[342]), .out(n344) );
  inv U1370 ( .a(b[343]), .out(n345) );
  inv U1371 ( .a(b[344]), .out(n346) );
  inv U1372 ( .a(b[345]), .out(n347) );
  inv U1373 ( .a(b[346]), .out(n348) );
  inv U1374 ( .a(b[347]), .out(n349) );
  inv U1375 ( .a(b[348]), .out(n350) );
  inv U1376 ( .a(b[349]), .out(n351) );
  inv U1377 ( .a(b[350]), .out(n352) );
  inv U1378 ( .a(b[351]), .out(n353) );
  inv U1379 ( .a(b[352]), .out(n354) );
  inv U1380 ( .a(b[353]), .out(n355) );
  inv U1381 ( .a(b[354]), .out(n356) );
  inv U1382 ( .a(b[355]), .out(n357) );
  inv U1383 ( .a(b[356]), .out(n358) );
  inv U1384 ( .a(b[357]), .out(n359) );
  inv U1385 ( .a(b[358]), .out(n360) );
  inv U1386 ( .a(b[359]), .out(n361) );
  inv U1387 ( .a(b[360]), .out(n362) );
  inv U1388 ( .a(b[361]), .out(n363) );
  inv U1389 ( .a(b[362]), .out(n364) );
  inv U1390 ( .a(b[363]), .out(n365) );
  inv U1391 ( .a(b[364]), .out(n366) );
  inv U1392 ( .a(b[365]), .out(n367) );
  inv U1393 ( .a(b[366]), .out(n368) );
  inv U1394 ( .a(b[367]), .out(n369) );
  inv U1395 ( .a(b[368]), .out(n370) );
  inv U1396 ( .a(b[369]), .out(n371) );
  inv U1397 ( .a(b[370]), .out(n372) );
  inv U1398 ( .a(b[371]), .out(n373) );
  inv U1399 ( .a(b[372]), .out(n374) );
  inv U1400 ( .a(b[373]), .out(n375) );
  inv U1401 ( .a(b[374]), .out(n376) );
  inv U1402 ( .a(b[375]), .out(n377) );
  inv U1403 ( .a(b[376]), .out(n378) );
  inv U1404 ( .a(b[377]), .out(n379) );
  inv U1405 ( .a(b[378]), .out(n380) );
  inv U1406 ( .a(b[379]), .out(n381) );
  inv U1407 ( .a(b[380]), .out(n382) );
  inv U1408 ( .a(b[381]), .out(n383) );
  inv U1409 ( .a(b[382]), .out(n384) );
  inv U1410 ( .a(b[383]), .out(n385) );
  inv U1411 ( .a(b[384]), .out(n386) );
  inv U1412 ( .a(b[385]), .out(n387) );
  inv U1413 ( .a(b[386]), .out(n388) );
  inv U1414 ( .a(b[387]), .out(n389) );
  inv U1415 ( .a(b[388]), .out(n390) );
  inv U1416 ( .a(b[389]), .out(n391) );
  inv U1417 ( .a(b[390]), .out(n392) );
  inv U1418 ( .a(b[391]), .out(n393) );
  inv U1419 ( .a(b[392]), .out(n394) );
  inv U1420 ( .a(b[393]), .out(n395) );
  inv U1421 ( .a(b[394]), .out(n396) );
  inv U1422 ( .a(b[395]), .out(n397) );
  inv U1423 ( .a(b[396]), .out(n398) );
  inv U1424 ( .a(b[397]), .out(n399) );
  inv U1425 ( .a(b[398]), .out(n400) );
  inv U1426 ( .a(b[399]), .out(n401) );
  inv U1427 ( .a(b[400]), .out(n402) );
  inv U1428 ( .a(b[401]), .out(n403) );
  inv U1429 ( .a(b[402]), .out(n404) );
  inv U1430 ( .a(b[403]), .out(n405) );
  inv U1431 ( .a(b[404]), .out(n406) );
  inv U1432 ( .a(b[405]), .out(n407) );
  inv U1433 ( .a(b[406]), .out(n408) );
  inv U1434 ( .a(b[407]), .out(n409) );
  inv U1435 ( .a(b[408]), .out(n410) );
  inv U1436 ( .a(b[409]), .out(n411) );
  inv U1437 ( .a(b[410]), .out(n412) );
  inv U1438 ( .a(b[411]), .out(n413) );
  inv U1439 ( .a(b[412]), .out(n414) );
  inv U1440 ( .a(b[413]), .out(n415) );
  inv U1441 ( .a(b[414]), .out(n416) );
  inv U1442 ( .a(b[415]), .out(n417) );
  inv U1443 ( .a(b[416]), .out(n418) );
  inv U1444 ( .a(b[417]), .out(n419) );
  inv U1445 ( .a(b[418]), .out(n420) );
  inv U1446 ( .a(b[419]), .out(n421) );
  inv U1447 ( .a(b[420]), .out(n422) );
  inv U1448 ( .a(b[421]), .out(n423) );
  inv U1449 ( .a(b[422]), .out(n424) );
  inv U1450 ( .a(b[423]), .out(n425) );
  inv U1451 ( .a(b[424]), .out(n426) );
  inv U1452 ( .a(b[425]), .out(n427) );
  inv U1453 ( .a(b[426]), .out(n428) );
  inv U1454 ( .a(b[427]), .out(n429) );
  inv U1455 ( .a(b[428]), .out(n430) );
  inv U1456 ( .a(b[429]), .out(n431) );
  inv U1457 ( .a(b[430]), .out(n432) );
  inv U1458 ( .a(b[431]), .out(n433) );
  inv U1459 ( .a(b[432]), .out(n434) );
  inv U1460 ( .a(b[433]), .out(n435) );
  inv U1461 ( .a(b[434]), .out(n436) );
  inv U1462 ( .a(b[435]), .out(n437) );
  inv U1463 ( .a(b[436]), .out(n438) );
  inv U1464 ( .a(b[437]), .out(n439) );
  inv U1465 ( .a(b[438]), .out(n440) );
  inv U1466 ( .a(b[439]), .out(n441) );
  inv U1467 ( .a(b[440]), .out(n442) );
  inv U1468 ( .a(b[441]), .out(n443) );
  inv U1469 ( .a(b[442]), .out(n444) );
  inv U1470 ( .a(b[443]), .out(n445) );
  inv U1471 ( .a(b[444]), .out(n446) );
  inv U1472 ( .a(b[445]), .out(n447) );
  inv U1473 ( .a(b[446]), .out(n448) );
  inv U1474 ( .a(b[447]), .out(n449) );
  inv U1475 ( .a(b[448]), .out(n450) );
  inv U1476 ( .a(b[449]), .out(n451) );
  inv U1477 ( .a(b[450]), .out(n452) );
  inv U1478 ( .a(b[451]), .out(n453) );
  inv U1479 ( .a(b[452]), .out(n454) );
  inv U1480 ( .a(b[453]), .out(n455) );
  inv U1481 ( .a(b[454]), .out(n456) );
  inv U1482 ( .a(b[455]), .out(n457) );
  inv U1483 ( .a(b[456]), .out(n458) );
  inv U1484 ( .a(b[457]), .out(n459) );
  inv U1485 ( .a(b[458]), .out(n460) );
  inv U1486 ( .a(b[459]), .out(n461) );
  inv U1487 ( .a(b[460]), .out(n462) );
  inv U1488 ( .a(b[461]), .out(n463) );
  inv U1489 ( .a(b[462]), .out(n464) );
  inv U1490 ( .a(b[463]), .out(n465) );
  inv U1491 ( .a(b[464]), .out(n466) );
  inv U1492 ( .a(b[465]), .out(n467) );
  inv U1493 ( .a(b[466]), .out(n468) );
  inv U1494 ( .a(b[467]), .out(n469) );
  inv U1495 ( .a(b[468]), .out(n470) );
  inv U1496 ( .a(b[469]), .out(n471) );
  inv U1497 ( .a(b[470]), .out(n472) );
  inv U1498 ( .a(b[471]), .out(n473) );
  inv U1499 ( .a(b[472]), .out(n474) );
  inv U1500 ( .a(b[473]), .out(n475) );
  inv U1501 ( .a(b[474]), .out(n476) );
  inv U1502 ( .a(b[475]), .out(n477) );
  inv U1503 ( .a(b[476]), .out(n478) );
  inv U1504 ( .a(b[477]), .out(n479) );
  inv U1505 ( .a(b[478]), .out(n480) );
  inv U1506 ( .a(b[479]), .out(n481) );
  inv U1507 ( .a(b[480]), .out(n482) );
  inv U1508 ( .a(b[481]), .out(n483) );
  inv U1509 ( .a(b[482]), .out(n484) );
  inv U1510 ( .a(b[483]), .out(n485) );
  inv U1511 ( .a(b[484]), .out(n486) );
  inv U1512 ( .a(b[485]), .out(n487) );
  inv U1513 ( .a(b[486]), .out(n488) );
  inv U1514 ( .a(b[487]), .out(n489) );
  inv U1515 ( .a(b[488]), .out(n490) );
  inv U1516 ( .a(b[489]), .out(n491) );
  inv U1517 ( .a(b[490]), .out(n492) );
  inv U1518 ( .a(b[491]), .out(n493) );
  inv U1519 ( .a(b[492]), .out(n494) );
  inv U1520 ( .a(b[493]), .out(n495) );
  inv U1521 ( .a(b[494]), .out(n496) );
  inv U1522 ( .a(b[495]), .out(n497) );
  inv U1523 ( .a(b[496]), .out(n498) );
  inv U1524 ( .a(b[497]), .out(n499) );
  inv U1525 ( .a(b[498]), .out(n500) );
  inv U1526 ( .a(b[499]), .out(n501) );
  inv U1527 ( .a(b[500]), .out(n502) );
  inv U1528 ( .a(b[501]), .out(n503) );
  inv U1529 ( .a(b[502]), .out(n504) );
  inv U1530 ( .a(b[503]), .out(n505) );
  inv U1531 ( .a(b[504]), .out(n506) );
  inv U1532 ( .a(b[505]), .out(n507) );
  inv U1533 ( .a(b[506]), .out(n508) );
  inv U1534 ( .a(b[507]), .out(n509) );
  inv U1535 ( .a(b[508]), .out(n510) );
  inv U1536 ( .a(b[509]), .out(n511) );
  inv U1537 ( .a(b[510]), .out(n512) );
  inv U1538 ( .a(b[511]), .out(n513) );
  inv U1539 ( .a(b[512]), .out(n514) );
  inv U1540 ( .a(b[513]), .out(n515) );
  inv U1541 ( .a(b[514]), .out(n516) );
  inv U1542 ( .a(b[515]), .out(n517) );
  inv U1543 ( .a(b[516]), .out(n518) );
  inv U1544 ( .a(b[517]), .out(n519) );
  inv U1545 ( .a(b[518]), .out(n520) );
  inv U1546 ( .a(b[519]), .out(n521) );
  inv U1547 ( .a(b[520]), .out(n522) );
  inv U1548 ( .a(b[521]), .out(n523) );
  inv U1549 ( .a(b[522]), .out(n524) );
  inv U1550 ( .a(b[523]), .out(n525) );
  inv U1551 ( .a(b[524]), .out(n526) );
  inv U1552 ( .a(b[525]), .out(n527) );
  inv U1553 ( .a(b[526]), .out(n528) );
  inv U1554 ( .a(b[527]), .out(n529) );
  inv U1555 ( .a(b[528]), .out(n530) );
  inv U1556 ( .a(b[529]), .out(n531) );
  inv U1557 ( .a(b[530]), .out(n532) );
  inv U1558 ( .a(b[531]), .out(n533) );
  inv U1559 ( .a(b[532]), .out(n534) );
  inv U1560 ( .a(b[533]), .out(n535) );
  inv U1561 ( .a(b[534]), .out(n536) );
  inv U1562 ( .a(b[535]), .out(n537) );
  inv U1563 ( .a(b[536]), .out(n538) );
  inv U1564 ( .a(b[537]), .out(n539) );
  inv U1565 ( .a(b[538]), .out(n540) );
  inv U1566 ( .a(b[539]), .out(n541) );
  inv U1567 ( .a(b[540]), .out(n542) );
  inv U1568 ( .a(b[541]), .out(n543) );
  inv U1569 ( .a(b[542]), .out(n544) );
  inv U1570 ( .a(b[543]), .out(n545) );
  inv U1571 ( .a(b[544]), .out(n546) );
  inv U1572 ( .a(b[545]), .out(n547) );
  inv U1573 ( .a(b[546]), .out(n548) );
  inv U1574 ( .a(b[547]), .out(n549) );
  inv U1575 ( .a(b[548]), .out(n550) );
  inv U1576 ( .a(b[549]), .out(n551) );
  inv U1577 ( .a(b[550]), .out(n552) );
  inv U1578 ( .a(b[551]), .out(n553) );
  inv U1579 ( .a(b[552]), .out(n554) );
  inv U1580 ( .a(b[553]), .out(n555) );
  inv U1581 ( .a(b[554]), .out(n556) );
  inv U1582 ( .a(b[555]), .out(n557) );
  inv U1583 ( .a(b[556]), .out(n558) );
  inv U1584 ( .a(b[557]), .out(n559) );
  inv U1585 ( .a(b[558]), .out(n560) );
  inv U1586 ( .a(b[559]), .out(n561) );
  inv U1587 ( .a(b[560]), .out(n562) );
  inv U1588 ( .a(b[561]), .out(n563) );
  inv U1589 ( .a(b[562]), .out(n564) );
  inv U1590 ( .a(b[563]), .out(n565) );
  inv U1591 ( .a(b[564]), .out(n566) );
  inv U1592 ( .a(b[565]), .out(n567) );
  inv U1593 ( .a(b[566]), .out(n568) );
  inv U1594 ( .a(b[567]), .out(n569) );
  inv U1595 ( .a(b[568]), .out(n570) );
  inv U1596 ( .a(b[569]), .out(n571) );
  inv U1597 ( .a(b[570]), .out(n572) );
  inv U1598 ( .a(b[571]), .out(n573) );
  inv U1599 ( .a(b[572]), .out(n574) );
  inv U1600 ( .a(b[573]), .out(n575) );
  inv U1601 ( .a(b[574]), .out(n576) );
  inv U1602 ( .a(b[575]), .out(n577) );
  inv U1603 ( .a(b[576]), .out(n578) );
  inv U1604 ( .a(b[577]), .out(n579) );
  inv U1605 ( .a(b[578]), .out(n580) );
  inv U1606 ( .a(b[579]), .out(n581) );
  inv U1607 ( .a(b[580]), .out(n582) );
  inv U1608 ( .a(b[581]), .out(n583) );
  inv U1609 ( .a(b[582]), .out(n584) );
  inv U1610 ( .a(b[583]), .out(n585) );
  inv U1611 ( .a(b[584]), .out(n586) );
  inv U1612 ( .a(b[585]), .out(n587) );
  inv U1613 ( .a(b[586]), .out(n588) );
  inv U1614 ( .a(b[587]), .out(n589) );
  inv U1615 ( .a(b[588]), .out(n590) );
  inv U1616 ( .a(b[589]), .out(n591) );
  inv U1617 ( .a(b[590]), .out(n592) );
  inv U1618 ( .a(b[591]), .out(n593) );
  inv U1619 ( .a(b[592]), .out(n594) );
  inv U1620 ( .a(b[593]), .out(n595) );
  inv U1621 ( .a(b[594]), .out(n596) );
  inv U1622 ( .a(b[595]), .out(n597) );
  inv U1623 ( .a(b[596]), .out(n598) );
  inv U1624 ( .a(b[597]), .out(n599) );
  inv U1625 ( .a(b[598]), .out(n600) );
  inv U1626 ( .a(b[599]), .out(n601) );
  inv U1627 ( .a(b[600]), .out(n602) );
  inv U1628 ( .a(b[601]), .out(n603) );
  inv U1629 ( .a(b[602]), .out(n604) );
  inv U1630 ( .a(b[603]), .out(n605) );
  inv U1631 ( .a(b[604]), .out(n606) );
  inv U1632 ( .a(b[605]), .out(n607) );
  inv U1633 ( .a(b[606]), .out(n608) );
  inv U1634 ( .a(b[607]), .out(n609) );
  inv U1635 ( .a(b[608]), .out(n610) );
  inv U1636 ( .a(b[609]), .out(n611) );
  inv U1637 ( .a(b[610]), .out(n612) );
  inv U1638 ( .a(b[611]), .out(n613) );
  inv U1639 ( .a(b[612]), .out(n614) );
  inv U1640 ( .a(b[613]), .out(n615) );
  inv U1641 ( .a(b[614]), .out(n616) );
  inv U1642 ( .a(b[615]), .out(n617) );
  inv U1643 ( .a(b[616]), .out(n618) );
  inv U1644 ( .a(b[617]), .out(n619) );
  inv U1645 ( .a(b[618]), .out(n620) );
  inv U1646 ( .a(b[619]), .out(n621) );
  inv U1647 ( .a(b[620]), .out(n622) );
  inv U1648 ( .a(b[621]), .out(n623) );
  inv U1649 ( .a(b[622]), .out(n624) );
  inv U1650 ( .a(b[623]), .out(n625) );
  inv U1651 ( .a(b[624]), .out(n626) );
  inv U1652 ( .a(b[625]), .out(n627) );
  inv U1653 ( .a(b[626]), .out(n628) );
  inv U1654 ( .a(b[627]), .out(n629) );
  inv U1655 ( .a(b[628]), .out(n630) );
  inv U1656 ( .a(b[629]), .out(n631) );
  inv U1657 ( .a(b[630]), .out(n632) );
  inv U1658 ( .a(b[631]), .out(n633) );
  inv U1659 ( .a(b[632]), .out(n634) );
  inv U1660 ( .a(b[633]), .out(n635) );
  inv U1661 ( .a(b[634]), .out(n636) );
  inv U1662 ( .a(b[635]), .out(n637) );
  inv U1663 ( .a(b[636]), .out(n638) );
  inv U1664 ( .a(b[637]), .out(n639) );
  inv U1665 ( .a(b[638]), .out(n640) );
  inv U1666 ( .a(b[639]), .out(n641) );
  inv U1667 ( .a(b[640]), .out(n642) );
  inv U1668 ( .a(b[641]), .out(n643) );
  inv U1669 ( .a(b[642]), .out(n644) );
  inv U1670 ( .a(b[643]), .out(n645) );
  inv U1671 ( .a(b[644]), .out(n646) );
  inv U1672 ( .a(b[645]), .out(n647) );
  inv U1673 ( .a(b[646]), .out(n648) );
  inv U1674 ( .a(b[647]), .out(n649) );
  inv U1675 ( .a(b[648]), .out(n650) );
  inv U1676 ( .a(b[649]), .out(n651) );
  inv U1677 ( .a(b[650]), .out(n652) );
  inv U1678 ( .a(b[651]), .out(n653) );
  inv U1679 ( .a(b[652]), .out(n654) );
  inv U1680 ( .a(b[653]), .out(n655) );
  inv U1681 ( .a(b[654]), .out(n656) );
  inv U1682 ( .a(b[655]), .out(n657) );
  inv U1683 ( .a(b[656]), .out(n658) );
  inv U1684 ( .a(b[657]), .out(n659) );
  inv U1685 ( .a(b[658]), .out(n660) );
  inv U1686 ( .a(b[659]), .out(n661) );
  inv U1687 ( .a(b[660]), .out(n662) );
  inv U1688 ( .a(b[661]), .out(n663) );
  inv U1689 ( .a(b[662]), .out(n664) );
  inv U1690 ( .a(b[663]), .out(n665) );
  inv U1691 ( .a(b[664]), .out(n666) );
  inv U1692 ( .a(b[665]), .out(n667) );
  inv U1693 ( .a(b[666]), .out(n668) );
  inv U1694 ( .a(b[667]), .out(n669) );
  inv U1695 ( .a(b[668]), .out(n670) );
  inv U1696 ( .a(b[669]), .out(n671) );
  inv U1697 ( .a(b[670]), .out(n672) );
  inv U1698 ( .a(b[671]), .out(n673) );
  inv U1699 ( .a(b[672]), .out(n674) );
  inv U1700 ( .a(b[673]), .out(n675) );
  inv U1701 ( .a(b[674]), .out(n676) );
  inv U1702 ( .a(b[675]), .out(n677) );
  inv U1703 ( .a(b[676]), .out(n678) );
  inv U1704 ( .a(b[677]), .out(n679) );
  inv U1705 ( .a(b[678]), .out(n680) );
  inv U1706 ( .a(b[679]), .out(n681) );
  inv U1707 ( .a(b[680]), .out(n682) );
  inv U1708 ( .a(b[681]), .out(n683) );
  inv U1709 ( .a(b[682]), .out(n684) );
  inv U1710 ( .a(b[683]), .out(n685) );
  inv U1711 ( .a(b[684]), .out(n686) );
  inv U1712 ( .a(b[685]), .out(n687) );
  inv U1713 ( .a(b[686]), .out(n688) );
  inv U1714 ( .a(b[687]), .out(n689) );
  inv U1715 ( .a(b[688]), .out(n690) );
  inv U1716 ( .a(b[689]), .out(n691) );
  inv U1717 ( .a(b[690]), .out(n692) );
  inv U1718 ( .a(b[691]), .out(n693) );
  inv U1719 ( .a(b[692]), .out(n694) );
  inv U1720 ( .a(b[693]), .out(n695) );
  inv U1721 ( .a(b[694]), .out(n696) );
  inv U1722 ( .a(b[695]), .out(n697) );
  inv U1723 ( .a(b[696]), .out(n698) );
  inv U1724 ( .a(b[697]), .out(n699) );
  inv U1725 ( .a(b[698]), .out(n700) );
  inv U1726 ( .a(b[699]), .out(n701) );
  inv U1727 ( .a(b[700]), .out(n702) );
  inv U1728 ( .a(b[701]), .out(n703) );
  inv U1729 ( .a(b[702]), .out(n704) );
  inv U1730 ( .a(b[703]), .out(n705) );
  inv U1731 ( .a(b[704]), .out(n706) );
  inv U1732 ( .a(b[705]), .out(n707) );
  inv U1733 ( .a(b[706]), .out(n708) );
  inv U1734 ( .a(b[707]), .out(n709) );
  inv U1735 ( .a(b[708]), .out(n710) );
  inv U1736 ( .a(b[709]), .out(n711) );
  inv U1737 ( .a(b[710]), .out(n712) );
  inv U1738 ( .a(b[711]), .out(n713) );
  inv U1739 ( .a(b[712]), .out(n714) );
  inv U1740 ( .a(b[713]), .out(n715) );
  inv U1741 ( .a(b[714]), .out(n716) );
  inv U1742 ( .a(b[715]), .out(n717) );
  inv U1743 ( .a(b[716]), .out(n718) );
  inv U1744 ( .a(b[717]), .out(n719) );
  inv U1745 ( .a(b[718]), .out(n720) );
  inv U1746 ( .a(b[719]), .out(n721) );
  inv U1747 ( .a(b[720]), .out(n722) );
  inv U1748 ( .a(b[721]), .out(n723) );
  inv U1749 ( .a(b[722]), .out(n724) );
  inv U1750 ( .a(b[723]), .out(n725) );
  inv U1751 ( .a(b[724]), .out(n726) );
  inv U1752 ( .a(b[725]), .out(n727) );
  inv U1753 ( .a(b[726]), .out(n728) );
  inv U1754 ( .a(b[727]), .out(n729) );
  inv U1755 ( .a(b[728]), .out(n730) );
  inv U1756 ( .a(b[729]), .out(n731) );
  inv U1757 ( .a(b[730]), .out(n732) );
  inv U1758 ( .a(b[731]), .out(n733) );
  inv U1759 ( .a(b[732]), .out(n734) );
  inv U1760 ( .a(b[733]), .out(n735) );
  inv U1761 ( .a(b[734]), .out(n736) );
  inv U1762 ( .a(b[735]), .out(n737) );
  inv U1763 ( .a(b[736]), .out(n738) );
  inv U1764 ( .a(b[737]), .out(n739) );
  inv U1765 ( .a(b[738]), .out(n740) );
  inv U1766 ( .a(b[739]), .out(n741) );
  inv U1767 ( .a(b[740]), .out(n742) );
  inv U1768 ( .a(b[741]), .out(n743) );
  inv U1769 ( .a(b[742]), .out(n744) );
  inv U1770 ( .a(b[743]), .out(n745) );
  inv U1771 ( .a(b[744]), .out(n746) );
  inv U1772 ( .a(b[745]), .out(n747) );
  inv U1773 ( .a(b[746]), .out(n748) );
  inv U1774 ( .a(b[747]), .out(n749) );
  inv U1775 ( .a(b[748]), .out(n750) );
  inv U1776 ( .a(b[749]), .out(n751) );
  inv U1777 ( .a(b[750]), .out(n752) );
  inv U1778 ( .a(b[751]), .out(n753) );
  inv U1779 ( .a(b[752]), .out(n754) );
  inv U1780 ( .a(b[753]), .out(n755) );
  inv U1781 ( .a(b[754]), .out(n756) );
  inv U1782 ( .a(b[755]), .out(n757) );
  inv U1783 ( .a(b[756]), .out(n758) );
  inv U1784 ( .a(b[757]), .out(n759) );
  inv U1785 ( .a(b[758]), .out(n760) );
  inv U1786 ( .a(b[759]), .out(n761) );
  inv U1787 ( .a(b[760]), .out(n762) );
  inv U1788 ( .a(b[761]), .out(n763) );
  inv U1789 ( .a(b[762]), .out(n764) );
  inv U1790 ( .a(b[763]), .out(n765) );
  inv U1791 ( .a(b[764]), .out(n766) );
  inv U1792 ( .a(b[765]), .out(n767) );
  inv U1793 ( .a(b[766]), .out(n768) );
  inv U1794 ( .a(b[767]), .out(n769) );
  inv U1795 ( .a(b[768]), .out(n770) );
  inv U1796 ( .a(b[769]), .out(n771) );
  inv U1797 ( .a(b[770]), .out(n772) );
  inv U1798 ( .a(b[771]), .out(n773) );
  inv U1799 ( .a(b[772]), .out(n774) );
  inv U1800 ( .a(b[773]), .out(n775) );
  inv U1801 ( .a(b[774]), .out(n776) );
  inv U1802 ( .a(b[775]), .out(n777) );
  inv U1803 ( .a(b[776]), .out(n778) );
  inv U1804 ( .a(b[777]), .out(n779) );
  inv U1805 ( .a(b[778]), .out(n780) );
  inv U1806 ( .a(b[779]), .out(n781) );
  inv U1807 ( .a(b[780]), .out(n782) );
  inv U1808 ( .a(b[781]), .out(n783) );
  inv U1809 ( .a(b[782]), .out(n784) );
  inv U1810 ( .a(b[783]), .out(n785) );
  inv U1811 ( .a(b[784]), .out(n786) );
  inv U1812 ( .a(b[785]), .out(n787) );
  inv U1813 ( .a(b[786]), .out(n788) );
  inv U1814 ( .a(b[787]), .out(n789) );
  inv U1815 ( .a(b[788]), .out(n790) );
  inv U1816 ( .a(b[789]), .out(n791) );
  inv U1817 ( .a(b[790]), .out(n792) );
  inv U1818 ( .a(b[791]), .out(n793) );
  inv U1819 ( .a(b[792]), .out(n794) );
  inv U1820 ( .a(b[793]), .out(n795) );
  inv U1821 ( .a(b[794]), .out(n796) );
  inv U1822 ( .a(b[795]), .out(n797) );
  inv U1823 ( .a(b[796]), .out(n798) );
  inv U1824 ( .a(b[797]), .out(n799) );
  inv U1825 ( .a(b[798]), .out(n800) );
  inv U1826 ( .a(b[799]), .out(n801) );
  inv U1827 ( .a(b[800]), .out(n802) );
  inv U1828 ( .a(b[801]), .out(n803) );
  inv U1829 ( .a(b[802]), .out(n804) );
  inv U1830 ( .a(b[803]), .out(n805) );
  inv U1831 ( .a(b[804]), .out(n806) );
  inv U1832 ( .a(b[805]), .out(n807) );
  inv U1833 ( .a(b[806]), .out(n808) );
  inv U1834 ( .a(b[807]), .out(n809) );
  inv U1835 ( .a(b[808]), .out(n810) );
  inv U1836 ( .a(b[809]), .out(n811) );
  inv U1837 ( .a(b[810]), .out(n812) );
  inv U1838 ( .a(b[811]), .out(n813) );
  inv U1839 ( .a(b[812]), .out(n814) );
  inv U1840 ( .a(b[813]), .out(n815) );
  inv U1841 ( .a(b[814]), .out(n816) );
  inv U1842 ( .a(b[815]), .out(n817) );
  inv U1843 ( .a(b[816]), .out(n818) );
  inv U1844 ( .a(b[817]), .out(n819) );
  inv U1845 ( .a(b[818]), .out(n820) );
  inv U1846 ( .a(b[819]), .out(n821) );
  inv U1847 ( .a(b[820]), .out(n822) );
  inv U1848 ( .a(b[821]), .out(n823) );
  inv U1849 ( .a(b[822]), .out(n824) );
  inv U1850 ( .a(b[823]), .out(n825) );
  inv U1851 ( .a(b[824]), .out(n826) );
  inv U1852 ( .a(b[825]), .out(n827) );
  inv U1853 ( .a(b[826]), .out(n828) );
  inv U1854 ( .a(b[827]), .out(n829) );
  inv U1855 ( .a(b[828]), .out(n830) );
  inv U1856 ( .a(b[829]), .out(n831) );
  inv U1857 ( .a(b[830]), .out(n832) );
  inv U1858 ( .a(b[831]), .out(n833) );
  inv U1859 ( .a(b[832]), .out(n834) );
  inv U1860 ( .a(b[833]), .out(n835) );
  inv U1861 ( .a(b[834]), .out(n836) );
  inv U1862 ( .a(b[835]), .out(n837) );
  inv U1863 ( .a(b[836]), .out(n838) );
  inv U1864 ( .a(b[837]), .out(n839) );
  inv U1865 ( .a(b[838]), .out(n840) );
  inv U1866 ( .a(b[839]), .out(n841) );
  inv U1867 ( .a(b[840]), .out(n842) );
  inv U1868 ( .a(b[841]), .out(n843) );
  inv U1869 ( .a(b[842]), .out(n844) );
  inv U1870 ( .a(b[843]), .out(n845) );
  inv U1871 ( .a(b[844]), .out(n846) );
  inv U1872 ( .a(b[845]), .out(n847) );
  inv U1873 ( .a(b[846]), .out(n848) );
  inv U1874 ( .a(b[847]), .out(n849) );
  inv U1875 ( .a(b[848]), .out(n850) );
  inv U1876 ( .a(b[849]), .out(n851) );
  inv U1877 ( .a(b[850]), .out(n852) );
  inv U1878 ( .a(b[851]), .out(n853) );
  inv U1879 ( .a(b[852]), .out(n854) );
  inv U1880 ( .a(b[853]), .out(n855) );
  inv U1881 ( .a(b[854]), .out(n856) );
  inv U1882 ( .a(b[855]), .out(n857) );
  inv U1883 ( .a(b[856]), .out(n858) );
  inv U1884 ( .a(b[857]), .out(n859) );
  inv U1885 ( .a(b[858]), .out(n860) );
  inv U1886 ( .a(b[859]), .out(n861) );
  inv U1887 ( .a(b[860]), .out(n862) );
  inv U1888 ( .a(b[861]), .out(n863) );
  inv U1889 ( .a(b[862]), .out(n864) );
  inv U1890 ( .a(b[863]), .out(n865) );
  inv U1891 ( .a(b[864]), .out(n866) );
  inv U1892 ( .a(b[865]), .out(n867) );
  inv U1893 ( .a(b[866]), .out(n868) );
  inv U1894 ( .a(b[867]), .out(n869) );
  inv U1895 ( .a(b[868]), .out(n870) );
  inv U1896 ( .a(b[869]), .out(n871) );
  inv U1897 ( .a(b[870]), .out(n872) );
  inv U1898 ( .a(b[871]), .out(n873) );
  inv U1899 ( .a(b[872]), .out(n874) );
  inv U1900 ( .a(b[873]), .out(n875) );
  inv U1901 ( .a(b[874]), .out(n876) );
  inv U1902 ( .a(b[875]), .out(n877) );
  inv U1903 ( .a(b[876]), .out(n878) );
  inv U1904 ( .a(b[877]), .out(n879) );
  inv U1905 ( .a(b[878]), .out(n880) );
  inv U1906 ( .a(b[879]), .out(n881) );
  inv U1907 ( .a(b[880]), .out(n882) );
  inv U1908 ( .a(b[881]), .out(n883) );
  inv U1909 ( .a(b[882]), .out(n884) );
  inv U1910 ( .a(b[883]), .out(n885) );
  inv U1911 ( .a(b[884]), .out(n886) );
  inv U1912 ( .a(b[885]), .out(n887) );
  inv U1913 ( .a(b[886]), .out(n888) );
  inv U1914 ( .a(b[887]), .out(n889) );
  inv U1915 ( .a(b[888]), .out(n890) );
  inv U1916 ( .a(b[889]), .out(n891) );
  inv U1917 ( .a(b[890]), .out(n892) );
  inv U1918 ( .a(b[891]), .out(n893) );
  inv U1919 ( .a(b[892]), .out(n894) );
  inv U1920 ( .a(b[893]), .out(n895) );
  inv U1921 ( .a(b[894]), .out(n896) );
  inv U1922 ( .a(b[895]), .out(n897) );
  inv U1923 ( .a(b[896]), .out(n898) );
  inv U1924 ( .a(b[897]), .out(n899) );
  inv U1925 ( .a(b[898]), .out(n900) );
  inv U1926 ( .a(b[899]), .out(n901) );
  inv U1927 ( .a(b[900]), .out(n902) );
  inv U1928 ( .a(b[901]), .out(n903) );
  inv U1929 ( .a(b[902]), .out(n904) );
  inv U1930 ( .a(b[903]), .out(n905) );
  inv U1931 ( .a(b[904]), .out(n906) );
  inv U1932 ( .a(b[905]), .out(n907) );
  inv U1933 ( .a(b[906]), .out(n908) );
  inv U1934 ( .a(b[907]), .out(n909) );
  inv U1935 ( .a(b[908]), .out(n910) );
  inv U1936 ( .a(b[909]), .out(n911) );
  inv U1937 ( .a(b[910]), .out(n912) );
  inv U1938 ( .a(b[911]), .out(n913) );
  inv U1939 ( .a(b[912]), .out(n914) );
  inv U1940 ( .a(b[913]), .out(n915) );
  inv U1941 ( .a(b[914]), .out(n916) );
  inv U1942 ( .a(b[915]), .out(n917) );
  inv U1943 ( .a(b[916]), .out(n918) );
  inv U1944 ( .a(b[917]), .out(n919) );
  inv U1945 ( .a(b[918]), .out(n920) );
  inv U1946 ( .a(b[919]), .out(n921) );
  inv U1947 ( .a(b[920]), .out(n922) );
  inv U1948 ( .a(b[921]), .out(n923) );
  inv U1949 ( .a(b[922]), .out(n924) );
  inv U1950 ( .a(b[923]), .out(n925) );
  inv U1951 ( .a(b[924]), .out(n926) );
  inv U1952 ( .a(b[925]), .out(n927) );
  inv U1953 ( .a(b[926]), .out(n928) );
  inv U1954 ( .a(b[927]), .out(n929) );
  inv U1955 ( .a(b[928]), .out(n930) );
  inv U1956 ( .a(b[929]), .out(n931) );
  inv U1957 ( .a(b[930]), .out(n932) );
  inv U1958 ( .a(b[931]), .out(n933) );
  inv U1959 ( .a(b[932]), .out(n934) );
  inv U1960 ( .a(b[933]), .out(n935) );
  inv U1961 ( .a(b[934]), .out(n936) );
  inv U1962 ( .a(b[935]), .out(n937) );
  inv U1963 ( .a(b[936]), .out(n938) );
  inv U1964 ( .a(b[937]), .out(n939) );
  inv U1965 ( .a(b[938]), .out(n940) );
  inv U1966 ( .a(b[939]), .out(n941) );
  inv U1967 ( .a(b[940]), .out(n942) );
  inv U1968 ( .a(b[941]), .out(n943) );
  inv U1969 ( .a(b[942]), .out(n944) );
  inv U1970 ( .a(b[943]), .out(n945) );
  inv U1971 ( .a(b[944]), .out(n946) );
  inv U1972 ( .a(b[945]), .out(n947) );
  inv U1973 ( .a(b[946]), .out(n948) );
  inv U1974 ( .a(b[947]), .out(n949) );
  inv U1975 ( .a(b[948]), .out(n950) );
  inv U1976 ( .a(b[949]), .out(n951) );
  inv U1977 ( .a(b[950]), .out(n952) );
  inv U1978 ( .a(b[951]), .out(n953) );
  inv U1979 ( .a(b[952]), .out(n954) );
  inv U1980 ( .a(b[953]), .out(n955) );
  inv U1981 ( .a(b[954]), .out(n956) );
  inv U1982 ( .a(b[955]), .out(n957) );
  inv U1983 ( .a(b[956]), .out(n958) );
  inv U1984 ( .a(b[957]), .out(n959) );
  inv U1985 ( .a(b[958]), .out(n960) );
  inv U1986 ( .a(b[959]), .out(n961) );
  inv U1987 ( .a(b[960]), .out(n962) );
  inv U1988 ( .a(b[961]), .out(n963) );
  inv U1989 ( .a(b[962]), .out(n964) );
  inv U1990 ( .a(b[963]), .out(n965) );
  inv U1991 ( .a(b[964]), .out(n966) );
  inv U1992 ( .a(b[965]), .out(n967) );
  inv U1993 ( .a(b[966]), .out(n968) );
  inv U1994 ( .a(b[967]), .out(n969) );
  inv U1995 ( .a(b[968]), .out(n970) );
  inv U1996 ( .a(b[969]), .out(n971) );
  inv U1997 ( .a(b[970]), .out(n972) );
  inv U1998 ( .a(b[971]), .out(n973) );
  inv U1999 ( .a(b[972]), .out(n974) );
  inv U2000 ( .a(b[973]), .out(n975) );
  inv U2001 ( .a(b[974]), .out(n976) );
  inv U2002 ( .a(b[975]), .out(n977) );
  inv U2003 ( .a(b[976]), .out(n978) );
  inv U2004 ( .a(b[977]), .out(n979) );
  inv U2005 ( .a(b[978]), .out(n980) );
  inv U2006 ( .a(b[979]), .out(n981) );
  inv U2007 ( .a(b[980]), .out(n982) );
  inv U2008 ( .a(b[981]), .out(n983) );
  inv U2009 ( .a(b[982]), .out(n984) );
  inv U2010 ( .a(b[983]), .out(n985) );
  inv U2011 ( .a(b[984]), .out(n986) );
  inv U2012 ( .a(b[985]), .out(n987) );
  inv U2013 ( .a(b[986]), .out(n988) );
  inv U2014 ( .a(b[987]), .out(n989) );
  inv U2015 ( .a(b[988]), .out(n990) );
  inv U2016 ( .a(b[989]), .out(n991) );
  inv U2017 ( .a(b[990]), .out(n992) );
  inv U2018 ( .a(b[991]), .out(n993) );
  inv U2019 ( .a(b[992]), .out(n994) );
  inv U2020 ( .a(b[993]), .out(n995) );
  inv U2021 ( .a(b[994]), .out(n996) );
  inv U2022 ( .a(b[995]), .out(n997) );
  inv U2023 ( .a(b[996]), .out(n998) );
  inv U2024 ( .a(b[997]), .out(n999) );
  inv U2025 ( .a(b[998]), .out(n1000) );
  inv U2026 ( .a(b[999]), .out(n1001) );
  inv U2027 ( .a(b[1000]), .out(n1002) );
  inv U2028 ( .a(b[1001]), .out(n1003) );
  inv U2029 ( .a(b[1002]), .out(n1004) );
  inv U2030 ( .a(b[1003]), .out(n1005) );
  inv U2031 ( .a(b[1004]), .out(n1006) );
  inv U2032 ( .a(b[1005]), .out(n1007) );
  inv U2033 ( .a(b[1006]), .out(n1008) );
  inv U2034 ( .a(b[1007]), .out(n1009) );
  inv U2035 ( .a(b[1008]), .out(n1010) );
  inv U2036 ( .a(b[1009]), .out(n1011) );
  inv U2037 ( .a(b[1010]), .out(n1012) );
  inv U2038 ( .a(b[1011]), .out(n1013) );
  inv U2039 ( .a(b[1012]), .out(n1014) );
  inv U2040 ( .a(b[1013]), .out(n1015) );
  inv U2041 ( .a(b[1014]), .out(n1016) );
  inv U2042 ( .a(b[1015]), .out(n1017) );
  inv U2043 ( .a(b[1016]), .out(n1018) );
  inv U2044 ( .a(b[1017]), .out(n1019) );
  inv U2045 ( .a(b[1018]), .out(n1020) );
  inv U2046 ( .a(b[1019]), .out(n1021) );
  inv U2047 ( .a(b[1020]), .out(n1022) );
  inv U2048 ( .a(b[1021]), .out(n1023) );
  inv U2049 ( .a(b[1022]), .out(n1024) );
endmodule

