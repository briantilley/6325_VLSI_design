$example HSPICE setup file

* transistor model and d_ff cell netlist
.include "~/cad/spice/model013.lib"
.include d_ff.sp

.global vdd! gnd!
.option post runlvl=5

.param vdd=1.2

* instantiate d flip-flop
uut D R clk Q d_ff

* voltage source
vdd vdd! gnd! 1.2v

* data
d-in D gnd! pwl(0ns 0 5ns 0 5.05ns vdd 25ns vdd 25.05ns 0
		41ns 0 41.05ns vdd 47 vdd 47.05ns 0 51ns 0 51.05ns vdd
		61ns vdd 61.05ns 0 67ns 0 67.05ns vdd 100ns vdd)

* reset
r-in R gnd! pwl(0ns vdd 2ns vdd 2.05ns 0 71ns 0 71.05ns vdd 100ns vdd)

* clock
c-in clk gnd! pulse(0 vdd 4.9ns 50ps 50ps 4.9ns 10ns)

* load capacitance
cout out gnd! 80f

* analysis
.tran 10ps 100ns

******************************** MEASUREMENTS ********************************

* t_su latching in 1
.measure tran t_su_1 trig v(D) val=vdd/2 cross=1 targ v(clk) val=vdd/2 cross=1

* t_su latching in 0
.measure tran t_su_0 trig v(D) val=vdd/2 cross=1 targ v(clk) val=vdd/2 cross=1

* t_hold latching in 1
.measure tran t_hld_1 trig v(D) val=vdd/2 cross=1 targ v(clk) val=vdd/2 cross=1

* t_hold latching in 0
.measure tran t_hld_0 trig v(D) val=vdd/2 cross=1 targ v(clk) val=vdd/2 cross=1

* t_clk->Q
.measure tran t_clk-Q trig v(clk) val=vdd/2 cross=1 targ v(Q) val=vdd/2 cross=1

* t_D
.measure t_d_0 param='t_su_0+t_clk-Q'
.measure t_d_1 param='t_su_1+t_clk-Q'

.end







* * 0ns 1.2v 1ns 1.2v 1.05ns 0v 6ns 0v 6.05ns 1.2v 12ns 1.2v

* * transient analysis
* .tr 100ps 12ns
* * example of parameter sweep, replace numeric value W of pfet with WP in invlvs.sp
* * .tr 100ps 12ns sweep WP 1u 9u 0.5u

* .measure tran trise trig v(in) val=0.6v fall=1 targ v(out) val=0.6v rise=1 $measure tlh at 0.6v
* .measure tran tfall trig v(in) val=0.6v rise=1 targ v(out) val=0.6v fall=1 $measure tpl at 0.6v
* .measure tavg param = '(trise+tfall)/2' $calculate average delay
* .measure tdiff param='abs(trise-tfall)' $calculate delay difference
* .measure delay param='max(trise,tfall)' $calculate worst case delay

* *  method 1
* .measure tran iavg avg i(vdd) from=0 to=10n $average current in one clock cycle
* .measure energy param='1.2*iavg*10n' $calculate energy in one clock cycle
* .measure edp1 param='abs(delay*energy)'

* *  method 2
* .measure tran t1 when v(in)=1.19 fall=1
* .measure tran t2 when v(out)=1.19 rise=1
* .measure tran t3 when v(in)=0.01 rise=1
* .measure tran t4 when v(out)=0.01 fall=1
* .measure tran i1 avg i(vdd) from=t1 to=t2 $average current when output rise
* .measure tran i2 avg i(vdd) from=t3 to=t4 $average current when output fall
* .measure energy1 param='1.2*i1*(t2-t1)' $calculate energy when output rise
* .measure energy2 param='1.2*i2*(t4-t3)' $calculate energy when output fall
* .measure energysum param='energy1+energy2'
* .measure edp2 param='abs(delay*energysum)'

* .end
